module SimpleLACore(
  input         clock,
  input         reset,
  input         io_ipi,
  input  [7:0]  io_interrupt,
  output        io_inst_req_valid,
  output [31:0] io_inst_req_bits_addr,
  input         io_inst_resp_valid,
  input  [31:0] io_inst_resp_bits,
  output        io_data_req_valid,
  output [3:0]  io_data_req_bits_wen,
  output [31:0] io_data_req_bits_addr,
  output [31:0] io_data_req_bits_wdata,
  output        io_data_req_bits_cacop,
  output        io_data_req_bits_preld,
  input         io_data_resp_valid,
  input  [31:0] io_data_resp_bits,
  output [31:0] io_debug_pc,
  output [3:0]  io_debug_wen,
  output [4:0]  io_debug_wnum,
  output [31:0] io_debug_wdata
);
  reg [31:0] GR [0:31];
  wire [31:0] GR_rj_MPORT_data;
  wire [4:0] GR_rj_MPORT_addr;
  wire [31:0] GR_rkd_MPORT_data;
  wire [4:0] GR_rkd_MPORT_addr;
  wire [31:0] GR_MPORT_data;
  wire [4:0] GR_MPORT_addr;
  wire  GR_MPORT_mask;
  wire  GR_MPORT_en;
  reg  idle;
  reg [31:0] PC;
  wire [31:0] PC4 = PC + 32'h4;
  reg [63:0] timer;
  wire [63:0] _timer_T_1 = timer + 64'h1;
  reg  iStallReg;
  reg  dStallReg;
  reg [1:0] crmd_DATM;
  reg [1:0] crmd_DATF;
  reg  crmd_PG;
  reg  crmd_DA;
  reg  crmd_IE;
  reg [1:0] crmd_PLV;
  reg  csrs_1_PIE;
  reg [1:0] csrs_1_PPLV;
  reg  csrs_2_FPE;
  reg [12:0] csrs_3_LIE;
  reg [8:0] csrs_4_EsubCode;
  reg [5:0] csrs_4_Ecode;
  reg  csrs_4_IS_0;
  reg  csrs_4_IS_1;
  reg  csrs_4_IS_2;
  reg  csrs_4_IS_3;
  reg  csrs_4_IS_4;
  reg  csrs_4_IS_5;
  reg  csrs_4_IS_6;
  reg  csrs_4_IS_7;
  reg  csrs_4_IS_8;
  reg  csrs_4_IS_9;
  reg  csrs_4_IS_11;
  reg  csrs_4_IS_12;
  reg [31:0] csrs_5_PC;
  reg [31:0] badv_VAddr;
  reg [25:0] csrs_7_VA;
  reg  csrs_8_NE;
  reg [5:0] csrs_8_PS;
  reg [4:0] csrs_8_Index;
  reg [18:0] csrs_9_VPPN;
  reg [23:0] csrs_10_PPN;
  reg  csrs_10_G;
  reg [1:0] csrs_10_MAT;
  reg [1:0] csrs_10_PLV;
  reg  csrs_10_D;
  reg  csrs_10_V;
  reg [23:0] csrs_11_PPN;
  reg  csrs_11_G;
  reg [1:0] csrs_11_MAT;
  reg [1:0] csrs_11_PLV;
  reg  csrs_11_D;
  reg  csrs_11_V;
  reg [9:0] asid_ASID;
  reg [19:0] csrs_13_Base;
  reg [19:0] csrs_14_Base;
  reg [31:0] csrs_17_Data;
  reg [31:0] csrs_18_Data;
  reg [31:0] csrs_19_Data;
  reg [31:0] csrs_20_Data;
  reg [31:0] csrs_21_TID;
  reg [29:0] csrs_22_InitVal;
  reg  csrs_22_Periodic;
  reg  csrs_22_En;
  reg [31:0] csrs_23_TimeVal;
  reg  csrs_25_KLO;
  reg  csrs_25_ROLLB;
  reg [25:0] csrs_26_PA;
  reg [2:0] csrs_27_VSEG;
  reg [2:0] csrs_27_PSEG;
  reg [1:0] csrs_27_MAT;
  reg  csrs_27_PLV3;
  reg  csrs_27_PLV0;
  reg [2:0] csrs_28_VSEG;
  reg [2:0] csrs_28_PSEG;
  reg [1:0] csrs_28_MAT;
  reg  csrs_28_PLV3;
  reg  csrs_28_PLV0;
  wire [31:0] _tval_TimeVal_T_1 = csrs_23_TimeVal - 32'h1;
  wire [31:0] _tval_TimeVal_T_2 = {csrs_22_InitVal,2'h0};
  wire [31:0] _GEN_0 = csrs_22_Periodic ? _tval_TimeVal_T_2 : csrs_23_TimeVal;
  wire  _GEN_1 = csrs_22_Periodic & csrs_22_En;
  wire [31:0] _GEN_2 = csrs_23_TimeVal != 32'h0 ? _tval_TimeVal_T_1 : _GEN_0;
  wire  _GEN_3 = csrs_23_TimeVal != 32'h0 ? csrs_4_IS_11 : 1'h1;
  wire  _GEN_4 = csrs_23_TimeVal != 32'h0 ? csrs_22_En : _GEN_1;
  wire [31:0] _GEN_5 = csrs_22_En ? _GEN_2 : csrs_23_TimeVal;
  wire  _GEN_6 = csrs_22_En ? _GEN_3 : csrs_4_IS_11;
  wire  _GEN_7 = csrs_22_En ? _GEN_4 : csrs_22_En;
  wire [5:0] hi_lo = {csrs_4_IS_5,csrs_4_IS_4,csrs_4_IS_3,csrs_4_IS_2,csrs_4_IS_1,csrs_4_IS_0};
  wire [12:0] _hi_T = {csrs_4_IS_12,csrs_4_IS_11,1'h0,csrs_4_IS_9,csrs_4_IS_8,csrs_4_IS_7,csrs_4_IS_6,hi_lo};
  wire [12:0] _hi_T_1 = csrs_3_LIE & _hi_T;
  wire  INT = |_hi_T_1 & crmd_IE;
  wire  _T_27 = ~idle;
  wire  _T_32 = crmd_PLV != 2'h0;
  wire  _T_34 = PC[1:0] != 2'h0 | PC[31] & crmd_PLV != 2'h0;
  wire  _T_11 = crmd_PLV == 2'h0;
  wire  _T_13 = crmd_PLV == 2'h3;
  reg  tlb_0_E;
  reg [18:0] tlb_0_VPPN;
  reg [5:0] tlb_0_PS;
  wire  vaMatch_0 = tlb_0_VPPN[18:10] == PC[31:23] & (tlb_0_PS == 6'h16 | tlb_0_VPPN[9:0] == PC[22:13]);
  reg  tlb_0_G;
  reg [9:0] tlb_0_ASID;
  wire  asidMatch_0 = tlb_0_ASID == asid_ASID;
  wire  tlbHit_0 = tlb_0_E & vaMatch_0 & (tlb_0_G | asidMatch_0);
  reg  tlb_1_E;
  reg [18:0] tlb_1_VPPN;
  reg [5:0] tlb_1_PS;
  wire  vaMatch_1 = tlb_1_VPPN[18:10] == PC[31:23] & (tlb_1_PS == 6'h16 | tlb_1_VPPN[9:0] == PC[22:13]);
  reg  tlb_1_G;
  reg [9:0] tlb_1_ASID;
  wire  asidMatch_1 = tlb_1_ASID == asid_ASID;
  wire  tlbHit_1 = tlb_1_E & vaMatch_1 & (tlb_1_G | asidMatch_1);
  reg  tlb_2_E;
  reg [18:0] tlb_2_VPPN;
  reg [5:0] tlb_2_PS;
  wire  vaMatch_2 = tlb_2_VPPN[18:10] == PC[31:23] & (tlb_2_PS == 6'h16 | tlb_2_VPPN[9:0] == PC[22:13]);
  reg  tlb_2_G;
  reg [9:0] tlb_2_ASID;
  wire  asidMatch_2 = tlb_2_ASID == asid_ASID;
  wire  tlbHit_2 = tlb_2_E & vaMatch_2 & (tlb_2_G | asidMatch_2);
  reg  tlb_3_E;
  reg [18:0] tlb_3_VPPN;
  reg [5:0] tlb_3_PS;
  wire  vaMatch_3 = tlb_3_VPPN[18:10] == PC[31:23] & (tlb_3_PS == 6'h16 | tlb_3_VPPN[9:0] == PC[22:13]);
  reg  tlb_3_G;
  reg [9:0] tlb_3_ASID;
  wire  asidMatch_3 = tlb_3_ASID == asid_ASID;
  wire  tlbHit_3 = tlb_3_E & vaMatch_3 & (tlb_3_G | asidMatch_3);
  reg  tlb_4_E;
  reg [18:0] tlb_4_VPPN;
  reg [5:0] tlb_4_PS;
  wire  vaMatch_4 = tlb_4_VPPN[18:10] == PC[31:23] & (tlb_4_PS == 6'h16 | tlb_4_VPPN[9:0] == PC[22:13]);
  reg  tlb_4_G;
  reg [9:0] tlb_4_ASID;
  wire  asidMatch_4 = tlb_4_ASID == asid_ASID;
  wire  tlbHit_4 = tlb_4_E & vaMatch_4 & (tlb_4_G | asidMatch_4);
  reg  tlb_5_E;
  reg [18:0] tlb_5_VPPN;
  reg [5:0] tlb_5_PS;
  wire  vaMatch_5 = tlb_5_VPPN[18:10] == PC[31:23] & (tlb_5_PS == 6'h16 | tlb_5_VPPN[9:0] == PC[22:13]);
  reg  tlb_5_G;
  reg [9:0] tlb_5_ASID;
  wire  asidMatch_5 = tlb_5_ASID == asid_ASID;
  wire  tlbHit_5 = tlb_5_E & vaMatch_5 & (tlb_5_G | asidMatch_5);
  reg  tlb_6_E;
  reg [18:0] tlb_6_VPPN;
  reg [5:0] tlb_6_PS;
  wire  vaMatch_6 = tlb_6_VPPN[18:10] == PC[31:23] & (tlb_6_PS == 6'h16 | tlb_6_VPPN[9:0] == PC[22:13]);
  reg  tlb_6_G;
  reg [9:0] tlb_6_ASID;
  wire  asidMatch_6 = tlb_6_ASID == asid_ASID;
  wire  tlbHit_6 = tlb_6_E & vaMatch_6 & (tlb_6_G | asidMatch_6);
  reg  tlb_7_E;
  reg [18:0] tlb_7_VPPN;
  reg [5:0] tlb_7_PS;
  wire  vaMatch_7 = tlb_7_VPPN[18:10] == PC[31:23] & (tlb_7_PS == 6'h16 | tlb_7_VPPN[9:0] == PC[22:13]);
  reg  tlb_7_G;
  reg [9:0] tlb_7_ASID;
  wire  asidMatch_7 = tlb_7_ASID == asid_ASID;
  wire  tlbHit_7 = tlb_7_E & vaMatch_7 & (tlb_7_G | asidMatch_7);
  reg  tlb_8_E;
  reg [18:0] tlb_8_VPPN;
  reg [5:0] tlb_8_PS;
  wire  vaMatch_8 = tlb_8_VPPN[18:10] == PC[31:23] & (tlb_8_PS == 6'h16 | tlb_8_VPPN[9:0] == PC[22:13]);
  reg  tlb_8_G;
  reg [9:0] tlb_8_ASID;
  wire  asidMatch_8 = tlb_8_ASID == asid_ASID;
  wire  tlbHit_8 = tlb_8_E & vaMatch_8 & (tlb_8_G | asidMatch_8);
  reg  tlb_9_E;
  reg [18:0] tlb_9_VPPN;
  reg [5:0] tlb_9_PS;
  wire  vaMatch_9 = tlb_9_VPPN[18:10] == PC[31:23] & (tlb_9_PS == 6'h16 | tlb_9_VPPN[9:0] == PC[22:13]);
  reg  tlb_9_G;
  reg [9:0] tlb_9_ASID;
  wire  asidMatch_9 = tlb_9_ASID == asid_ASID;
  wire  tlbHit_9 = tlb_9_E & vaMatch_9 & (tlb_9_G | asidMatch_9);
  reg  tlb_10_E;
  reg [18:0] tlb_10_VPPN;
  reg [5:0] tlb_10_PS;
  wire  vaMatch_10 = tlb_10_VPPN[18:10] == PC[31:23] & (tlb_10_PS == 6'h16 | tlb_10_VPPN[9:0] == PC[22:13]);
  reg  tlb_10_G;
  reg [9:0] tlb_10_ASID;
  wire  asidMatch_10 = tlb_10_ASID == asid_ASID;
  wire  tlbHit_10 = tlb_10_E & vaMatch_10 & (tlb_10_G | asidMatch_10);
  reg  tlb_11_E;
  reg [18:0] tlb_11_VPPN;
  reg [5:0] tlb_11_PS;
  wire  vaMatch_11 = tlb_11_VPPN[18:10] == PC[31:23] & (tlb_11_PS == 6'h16 | tlb_11_VPPN[9:0] == PC[22:13]);
  reg  tlb_11_G;
  reg [9:0] tlb_11_ASID;
  wire  asidMatch_11 = tlb_11_ASID == asid_ASID;
  wire  tlbHit_11 = tlb_11_E & vaMatch_11 & (tlb_11_G | asidMatch_11);
  reg  tlb_12_E;
  reg [18:0] tlb_12_VPPN;
  reg [5:0] tlb_12_PS;
  wire  vaMatch_12 = tlb_12_VPPN[18:10] == PC[31:23] & (tlb_12_PS == 6'h16 | tlb_12_VPPN[9:0] == PC[22:13]);
  reg  tlb_12_G;
  reg [9:0] tlb_12_ASID;
  wire  asidMatch_12 = tlb_12_ASID == asid_ASID;
  wire  tlbHit_12 = tlb_12_E & vaMatch_12 & (tlb_12_G | asidMatch_12);
  reg  tlb_13_E;
  reg [18:0] tlb_13_VPPN;
  reg [5:0] tlb_13_PS;
  wire  vaMatch_13 = tlb_13_VPPN[18:10] == PC[31:23] & (tlb_13_PS == 6'h16 | tlb_13_VPPN[9:0] == PC[22:13]);
  reg  tlb_13_G;
  reg [9:0] tlb_13_ASID;
  wire  asidMatch_13 = tlb_13_ASID == asid_ASID;
  wire  tlbHit_13 = tlb_13_E & vaMatch_13 & (tlb_13_G | asidMatch_13);
  reg  tlb_14_E;
  reg [18:0] tlb_14_VPPN;
  reg [5:0] tlb_14_PS;
  wire  vaMatch_14 = tlb_14_VPPN[18:10] == PC[31:23] & (tlb_14_PS == 6'h16 | tlb_14_VPPN[9:0] == PC[22:13]);
  reg  tlb_14_G;
  reg [9:0] tlb_14_ASID;
  wire  asidMatch_14 = tlb_14_ASID == asid_ASID;
  wire  tlbHit_14 = tlb_14_E & vaMatch_14 & (tlb_14_G | asidMatch_14);
  reg  tlb_15_E;
  reg [18:0] tlb_15_VPPN;
  reg [5:0] tlb_15_PS;
  wire  vaMatch_15 = tlb_15_VPPN[18:10] == PC[31:23] & (tlb_15_PS == 6'h16 | tlb_15_VPPN[9:0] == PC[22:13]);
  reg  tlb_15_G;
  reg [9:0] tlb_15_ASID;
  wire  asidMatch_15 = tlb_15_ASID == asid_ASID;
  wire  tlbHit_15 = tlb_15_E & vaMatch_15 & (tlb_15_G | asidMatch_15);
  reg  tlb_16_E;
  reg [18:0] tlb_16_VPPN;
  reg [5:0] tlb_16_PS;
  wire  vaMatch_16 = tlb_16_VPPN[18:10] == PC[31:23] & (tlb_16_PS == 6'h16 | tlb_16_VPPN[9:0] == PC[22:13]);
  reg  tlb_16_G;
  reg [9:0] tlb_16_ASID;
  wire  asidMatch_16 = tlb_16_ASID == asid_ASID;
  wire  tlbHit_16 = tlb_16_E & vaMatch_16 & (tlb_16_G | asidMatch_16);
  reg  tlb_17_E;
  reg [18:0] tlb_17_VPPN;
  reg [5:0] tlb_17_PS;
  wire  vaMatch_17 = tlb_17_VPPN[18:10] == PC[31:23] & (tlb_17_PS == 6'h16 | tlb_17_VPPN[9:0] == PC[22:13]);
  reg  tlb_17_G;
  reg [9:0] tlb_17_ASID;
  wire  asidMatch_17 = tlb_17_ASID == asid_ASID;
  wire  tlbHit_17 = tlb_17_E & vaMatch_17 & (tlb_17_G | asidMatch_17);
  reg  tlb_18_E;
  reg [18:0] tlb_18_VPPN;
  reg [5:0] tlb_18_PS;
  wire  vaMatch_18 = tlb_18_VPPN[18:10] == PC[31:23] & (tlb_18_PS == 6'h16 | tlb_18_VPPN[9:0] == PC[22:13]);
  reg  tlb_18_G;
  reg [9:0] tlb_18_ASID;
  wire  asidMatch_18 = tlb_18_ASID == asid_ASID;
  wire  tlbHit_18 = tlb_18_E & vaMatch_18 & (tlb_18_G | asidMatch_18);
  reg  tlb_19_E;
  reg [18:0] tlb_19_VPPN;
  reg [5:0] tlb_19_PS;
  wire  vaMatch_19 = tlb_19_VPPN[18:10] == PC[31:23] & (tlb_19_PS == 6'h16 | tlb_19_VPPN[9:0] == PC[22:13]);
  reg  tlb_19_G;
  reg [9:0] tlb_19_ASID;
  wire  asidMatch_19 = tlb_19_ASID == asid_ASID;
  wire  tlbHit_19 = tlb_19_E & vaMatch_19 & (tlb_19_G | asidMatch_19);
  reg  tlb_20_E;
  reg [18:0] tlb_20_VPPN;
  reg [5:0] tlb_20_PS;
  wire  vaMatch_20 = tlb_20_VPPN[18:10] == PC[31:23] & (tlb_20_PS == 6'h16 | tlb_20_VPPN[9:0] == PC[22:13]);
  reg  tlb_20_G;
  reg [9:0] tlb_20_ASID;
  wire  asidMatch_20 = tlb_20_ASID == asid_ASID;
  wire  tlbHit_20 = tlb_20_E & vaMatch_20 & (tlb_20_G | asidMatch_20);
  reg  tlb_21_E;
  reg [18:0] tlb_21_VPPN;
  reg [5:0] tlb_21_PS;
  wire  vaMatch_21 = tlb_21_VPPN[18:10] == PC[31:23] & (tlb_21_PS == 6'h16 | tlb_21_VPPN[9:0] == PC[22:13]);
  reg  tlb_21_G;
  reg [9:0] tlb_21_ASID;
  wire  asidMatch_21 = tlb_21_ASID == asid_ASID;
  wire  tlbHit_21 = tlb_21_E & vaMatch_21 & (tlb_21_G | asidMatch_21);
  reg  tlb_22_E;
  reg [18:0] tlb_22_VPPN;
  reg [5:0] tlb_22_PS;
  wire  vaMatch_22 = tlb_22_VPPN[18:10] == PC[31:23] & (tlb_22_PS == 6'h16 | tlb_22_VPPN[9:0] == PC[22:13]);
  reg  tlb_22_G;
  reg [9:0] tlb_22_ASID;
  wire  asidMatch_22 = tlb_22_ASID == asid_ASID;
  wire  tlbHit_22 = tlb_22_E & vaMatch_22 & (tlb_22_G | asidMatch_22);
  reg  tlb_23_E;
  reg [18:0] tlb_23_VPPN;
  reg [5:0] tlb_23_PS;
  wire  vaMatch_23 = tlb_23_VPPN[18:10] == PC[31:23] & (tlb_23_PS == 6'h16 | tlb_23_VPPN[9:0] == PC[22:13]);
  reg  tlb_23_G;
  reg [9:0] tlb_23_ASID;
  wire  asidMatch_23 = tlb_23_ASID == asid_ASID;
  wire  tlbHit_23 = tlb_23_E & vaMatch_23 & (tlb_23_G | asidMatch_23);
  reg  tlb_24_E;
  reg [18:0] tlb_24_VPPN;
  reg [5:0] tlb_24_PS;
  wire  vaMatch_24 = tlb_24_VPPN[18:10] == PC[31:23] & (tlb_24_PS == 6'h16 | tlb_24_VPPN[9:0] == PC[22:13]);
  reg  tlb_24_G;
  reg [9:0] tlb_24_ASID;
  wire  asidMatch_24 = tlb_24_ASID == asid_ASID;
  wire  tlbHit_24 = tlb_24_E & vaMatch_24 & (tlb_24_G | asidMatch_24);
  reg  tlb_25_E;
  reg [18:0] tlb_25_VPPN;
  reg [5:0] tlb_25_PS;
  wire  vaMatch_25 = tlb_25_VPPN[18:10] == PC[31:23] & (tlb_25_PS == 6'h16 | tlb_25_VPPN[9:0] == PC[22:13]);
  reg  tlb_25_G;
  reg [9:0] tlb_25_ASID;
  wire  asidMatch_25 = tlb_25_ASID == asid_ASID;
  wire  tlbHit_25 = tlb_25_E & vaMatch_25 & (tlb_25_G | asidMatch_25);
  reg  tlb_26_E;
  reg [18:0] tlb_26_VPPN;
  reg [5:0] tlb_26_PS;
  wire  vaMatch_26 = tlb_26_VPPN[18:10] == PC[31:23] & (tlb_26_PS == 6'h16 | tlb_26_VPPN[9:0] == PC[22:13]);
  reg  tlb_26_G;
  reg [9:0] tlb_26_ASID;
  wire  asidMatch_26 = tlb_26_ASID == asid_ASID;
  wire  tlbHit_26 = tlb_26_E & vaMatch_26 & (tlb_26_G | asidMatch_26);
  reg  tlb_27_E;
  reg [18:0] tlb_27_VPPN;
  reg [5:0] tlb_27_PS;
  wire  vaMatch_27 = tlb_27_VPPN[18:10] == PC[31:23] & (tlb_27_PS == 6'h16 | tlb_27_VPPN[9:0] == PC[22:13]);
  reg  tlb_27_G;
  reg [9:0] tlb_27_ASID;
  wire  asidMatch_27 = tlb_27_ASID == asid_ASID;
  wire  tlbHit_27 = tlb_27_E & vaMatch_27 & (tlb_27_G | asidMatch_27);
  reg  tlb_28_E;
  reg [18:0] tlb_28_VPPN;
  reg [5:0] tlb_28_PS;
  wire  vaMatch_28 = tlb_28_VPPN[18:10] == PC[31:23] & (tlb_28_PS == 6'h16 | tlb_28_VPPN[9:0] == PC[22:13]);
  reg  tlb_28_G;
  reg [9:0] tlb_28_ASID;
  wire  asidMatch_28 = tlb_28_ASID == asid_ASID;
  wire  tlbHit_28 = tlb_28_E & vaMatch_28 & (tlb_28_G | asidMatch_28);
  reg  tlb_29_E;
  reg [18:0] tlb_29_VPPN;
  reg [5:0] tlb_29_PS;
  wire  vaMatch_29 = tlb_29_VPPN[18:10] == PC[31:23] & (tlb_29_PS == 6'h16 | tlb_29_VPPN[9:0] == PC[22:13]);
  reg  tlb_29_G;
  reg [9:0] tlb_29_ASID;
  wire  asidMatch_29 = tlb_29_ASID == asid_ASID;
  wire  tlbHit_29 = tlb_29_E & vaMatch_29 & (tlb_29_G | asidMatch_29);
  reg  tlb_30_E;
  reg [18:0] tlb_30_VPPN;
  reg [5:0] tlb_30_PS;
  wire  vaMatch_30 = tlb_30_VPPN[18:10] == PC[31:23] & (tlb_30_PS == 6'h16 | tlb_30_VPPN[9:0] == PC[22:13]);
  reg  tlb_30_G;
  reg [9:0] tlb_30_ASID;
  wire  asidMatch_30 = tlb_30_ASID == asid_ASID;
  wire  tlbHit_30 = tlb_30_E & vaMatch_30 & (tlb_30_G | asidMatch_30);
  wire  _miss_T_29 = tlbHit_0 | tlbHit_1 | tlbHit_2 | tlbHit_3 | tlbHit_4 | tlbHit_5 | tlbHit_6 | tlbHit_7 | tlbHit_8 |
    tlbHit_9 | tlbHit_10 | tlbHit_11 | tlbHit_12 | tlbHit_13 | tlbHit_14 | tlbHit_15 | tlbHit_16 | tlbHit_17 | tlbHit_18
     | tlbHit_19 | tlbHit_20 | tlbHit_21 | tlbHit_22 | tlbHit_23 | tlbHit_24 | tlbHit_25 | tlbHit_26 | tlbHit_27 |
    tlbHit_28 | tlbHit_29 | tlbHit_30;
  reg  tlb_31_E;
  reg [18:0] tlb_31_VPPN;
  reg [5:0] tlb_31_PS;
  wire  vaMatch_31 = tlb_31_VPPN[18:10] == PC[31:23] & (tlb_31_PS == 6'h16 | tlb_31_VPPN[9:0] == PC[22:13]);
  reg  tlb_31_G;
  reg [9:0] tlb_31_ASID;
  wire  asidMatch_31 = tlb_31_ASID == asid_ASID;
  wire  tlbHit_31 = tlb_31_E & vaMatch_31 & (tlb_31_G | asidMatch_31);
  wire  _GEN_10 = PC[31:29] == csrs_28_VSEG & (csrs_28_PLV0 & _T_11 | csrs_28_PLV3 & _T_13) ? 1'h0 : ~(_miss_T_29 |
    tlbHit_31);
  wire  miss = PC[31:29] == csrs_27_VSEG & (csrs_27_PLV0 & crmd_PLV == 2'h0 | csrs_27_PLV3 & crmd_PLV == 2'h3) ? 1'h0 :
    _GEN_10;
  wire  _GEN_30 = crmd_DA ? 1'h0 : miss;
  wire  _GEN_35 = PC[1:0] != 2'h0 | PC[31] & crmd_PLV != 2'h0 ? 1'h0 : _GEN_30;
  wire  _GEN_40 = ~INT & ~idle & _GEN_35;
  wire  _GEN_45 = dStallReg | iStallReg ? 1'h0 : _GEN_40;
  wire [5:0] _foundTLB_T_819 = tlbHit_0 ? tlb_0_PS : 6'h0;
  wire [5:0] _foundTLB_T_820 = tlbHit_1 ? tlb_1_PS : 6'h0;
  wire [5:0] _foundTLB_T_851 = _foundTLB_T_819 | _foundTLB_T_820;
  wire [5:0] _foundTLB_T_821 = tlbHit_2 ? tlb_2_PS : 6'h0;
  wire [5:0] _foundTLB_T_852 = _foundTLB_T_851 | _foundTLB_T_821;
  wire [5:0] _foundTLB_T_822 = tlbHit_3 ? tlb_3_PS : 6'h0;
  wire [5:0] _foundTLB_T_853 = _foundTLB_T_852 | _foundTLB_T_822;
  wire [5:0] _foundTLB_T_823 = tlbHit_4 ? tlb_4_PS : 6'h0;
  wire [5:0] _foundTLB_T_854 = _foundTLB_T_853 | _foundTLB_T_823;
  wire [5:0] _foundTLB_T_824 = tlbHit_5 ? tlb_5_PS : 6'h0;
  wire [5:0] _foundTLB_T_855 = _foundTLB_T_854 | _foundTLB_T_824;
  wire [5:0] _foundTLB_T_825 = tlbHit_6 ? tlb_6_PS : 6'h0;
  wire [5:0] _foundTLB_T_856 = _foundTLB_T_855 | _foundTLB_T_825;
  wire [5:0] _foundTLB_T_826 = tlbHit_7 ? tlb_7_PS : 6'h0;
  wire [5:0] _foundTLB_T_857 = _foundTLB_T_856 | _foundTLB_T_826;
  wire [5:0] _foundTLB_T_827 = tlbHit_8 ? tlb_8_PS : 6'h0;
  wire [5:0] _foundTLB_T_858 = _foundTLB_T_857 | _foundTLB_T_827;
  wire [5:0] _foundTLB_T_828 = tlbHit_9 ? tlb_9_PS : 6'h0;
  wire [5:0] _foundTLB_T_859 = _foundTLB_T_858 | _foundTLB_T_828;
  wire [5:0] _foundTLB_T_829 = tlbHit_10 ? tlb_10_PS : 6'h0;
  wire [5:0] _foundTLB_T_860 = _foundTLB_T_859 | _foundTLB_T_829;
  wire [5:0] _foundTLB_T_830 = tlbHit_11 ? tlb_11_PS : 6'h0;
  wire [5:0] _foundTLB_T_861 = _foundTLB_T_860 | _foundTLB_T_830;
  wire [5:0] _foundTLB_T_831 = tlbHit_12 ? tlb_12_PS : 6'h0;
  wire [5:0] _foundTLB_T_862 = _foundTLB_T_861 | _foundTLB_T_831;
  wire [5:0] _foundTLB_T_832 = tlbHit_13 ? tlb_13_PS : 6'h0;
  wire [5:0] _foundTLB_T_863 = _foundTLB_T_862 | _foundTLB_T_832;
  wire [5:0] _foundTLB_T_833 = tlbHit_14 ? tlb_14_PS : 6'h0;
  wire [5:0] _foundTLB_T_864 = _foundTLB_T_863 | _foundTLB_T_833;
  wire [5:0] _foundTLB_T_834 = tlbHit_15 ? tlb_15_PS : 6'h0;
  wire [5:0] _foundTLB_T_865 = _foundTLB_T_864 | _foundTLB_T_834;
  wire [5:0] _foundTLB_T_835 = tlbHit_16 ? tlb_16_PS : 6'h0;
  wire [5:0] _foundTLB_T_866 = _foundTLB_T_865 | _foundTLB_T_835;
  wire [5:0] _foundTLB_T_836 = tlbHit_17 ? tlb_17_PS : 6'h0;
  wire [5:0] _foundTLB_T_867 = _foundTLB_T_866 | _foundTLB_T_836;
  wire [5:0] _foundTLB_T_837 = tlbHit_18 ? tlb_18_PS : 6'h0;
  wire [5:0] _foundTLB_T_868 = _foundTLB_T_867 | _foundTLB_T_837;
  wire [5:0] _foundTLB_T_838 = tlbHit_19 ? tlb_19_PS : 6'h0;
  wire [5:0] _foundTLB_T_869 = _foundTLB_T_868 | _foundTLB_T_838;
  wire [5:0] _foundTLB_T_839 = tlbHit_20 ? tlb_20_PS : 6'h0;
  wire [5:0] _foundTLB_T_870 = _foundTLB_T_869 | _foundTLB_T_839;
  wire [5:0] _foundTLB_T_840 = tlbHit_21 ? tlb_21_PS : 6'h0;
  wire [5:0] _foundTLB_T_871 = _foundTLB_T_870 | _foundTLB_T_840;
  wire [5:0] _foundTLB_T_841 = tlbHit_22 ? tlb_22_PS : 6'h0;
  wire [5:0] _foundTLB_T_872 = _foundTLB_T_871 | _foundTLB_T_841;
  wire [5:0] _foundTLB_T_842 = tlbHit_23 ? tlb_23_PS : 6'h0;
  wire [5:0] _foundTLB_T_873 = _foundTLB_T_872 | _foundTLB_T_842;
  wire [5:0] _foundTLB_T_843 = tlbHit_24 ? tlb_24_PS : 6'h0;
  wire [5:0] _foundTLB_T_874 = _foundTLB_T_873 | _foundTLB_T_843;
  wire [5:0] _foundTLB_T_844 = tlbHit_25 ? tlb_25_PS : 6'h0;
  wire [5:0] _foundTLB_T_875 = _foundTLB_T_874 | _foundTLB_T_844;
  wire [5:0] _foundTLB_T_845 = tlbHit_26 ? tlb_26_PS : 6'h0;
  wire [5:0] _foundTLB_T_876 = _foundTLB_T_875 | _foundTLB_T_845;
  wire [5:0] _foundTLB_T_846 = tlbHit_27 ? tlb_27_PS : 6'h0;
  wire [5:0] _foundTLB_T_877 = _foundTLB_T_876 | _foundTLB_T_846;
  wire [5:0] _foundTLB_T_847 = tlbHit_28 ? tlb_28_PS : 6'h0;
  wire [5:0] _foundTLB_T_878 = _foundTLB_T_877 | _foundTLB_T_847;
  wire [5:0] _foundTLB_T_848 = tlbHit_29 ? tlb_29_PS : 6'h0;
  wire [5:0] _foundTLB_T_879 = _foundTLB_T_878 | _foundTLB_T_848;
  wire [5:0] _foundTLB_T_849 = tlbHit_30 ? tlb_30_PS : 6'h0;
  wire [5:0] _foundTLB_T_880 = _foundTLB_T_879 | _foundTLB_T_849;
  wire [5:0] _foundTLB_T_850 = tlbHit_31 ? tlb_31_PS : 6'h0;
  wire [5:0] foundTLB_PS = _foundTLB_T_880 | _foundTLB_T_850;
  wire  _oddPG_T = foundTLB_PS == 6'hc;
  wire  oddPG = foundTLB_PS == 6'hc ? PC[12] : PC[22];
  reg  tlb_0_P1_V;
  reg  tlb_1_P1_V;
  reg  tlb_2_P1_V;
  reg  tlb_3_P1_V;
  reg  tlb_4_P1_V;
  reg  tlb_5_P1_V;
  reg  tlb_6_P1_V;
  reg  tlb_7_P1_V;
  reg  tlb_8_P1_V;
  reg  tlb_9_P1_V;
  reg  tlb_10_P1_V;
  reg  tlb_11_P1_V;
  reg  tlb_12_P1_V;
  reg  tlb_13_P1_V;
  reg  tlb_14_P1_V;
  reg  tlb_15_P1_V;
  wire  _foundTLB_T_15 = tlbHit_15 & tlb_15_P1_V;
  wire  _foundTLB_T_46 = tlbHit_0 & tlb_0_P1_V | tlbHit_1 & tlb_1_P1_V | tlbHit_2 & tlb_2_P1_V | tlbHit_3 & tlb_3_P1_V
     | tlbHit_4 & tlb_4_P1_V | tlbHit_5 & tlb_5_P1_V | tlbHit_6 & tlb_6_P1_V | tlbHit_7 & tlb_7_P1_V | tlbHit_8 &
    tlb_8_P1_V | tlbHit_9 & tlb_9_P1_V | tlbHit_10 & tlb_10_P1_V | tlbHit_11 & tlb_11_P1_V | tlbHit_12 & tlb_12_P1_V |
    tlbHit_13 & tlb_13_P1_V | tlbHit_14 & tlb_14_P1_V | _foundTLB_T_15;
  reg  tlb_16_P1_V;
  reg  tlb_17_P1_V;
  reg  tlb_18_P1_V;
  reg  tlb_19_P1_V;
  reg  tlb_20_P1_V;
  reg  tlb_21_P1_V;
  reg  tlb_22_P1_V;
  reg  tlb_23_P1_V;
  reg  tlb_24_P1_V;
  reg  tlb_25_P1_V;
  reg  tlb_26_P1_V;
  reg  tlb_27_P1_V;
  reg  tlb_28_P1_V;
  reg  tlb_29_P1_V;
  reg  tlb_30_P1_V;
  wire  _foundTLB_T_61 = _foundTLB_T_46 | tlbHit_16 & tlb_16_P1_V | tlbHit_17 & tlb_17_P1_V | tlbHit_18 & tlb_18_P1_V |
    tlbHit_19 & tlb_19_P1_V | tlbHit_20 & tlb_20_P1_V | tlbHit_21 & tlb_21_P1_V | tlbHit_22 & tlb_22_P1_V | tlbHit_23 &
    tlb_23_P1_V | tlbHit_24 & tlb_24_P1_V | tlbHit_25 & tlb_25_P1_V | tlbHit_26 & tlb_26_P1_V | tlbHit_27 & tlb_27_P1_V
     | tlbHit_28 & tlb_28_P1_V | tlbHit_29 & tlb_29_P1_V | tlbHit_30 & tlb_30_P1_V;
  reg  tlb_31_P1_V;
  wire  foundTLB_P1_V = _foundTLB_T_61 | tlbHit_31 & tlb_31_P1_V;
  reg  tlb_0_P0_V;
  reg  tlb_1_P0_V;
  reg  tlb_2_P0_V;
  reg  tlb_3_P0_V;
  reg  tlb_4_P0_V;
  reg  tlb_5_P0_V;
  reg  tlb_6_P0_V;
  reg  tlb_7_P0_V;
  reg  tlb_8_P0_V;
  reg  tlb_9_P0_V;
  reg  tlb_10_P0_V;
  reg  tlb_11_P0_V;
  reg  tlb_12_P0_V;
  reg  tlb_13_P0_V;
  reg  tlb_14_P0_V;
  reg  tlb_15_P0_V;
  wire  _foundTLB_T_330 = tlbHit_15 & tlb_15_P0_V;
  wire  _foundTLB_T_361 = tlbHit_0 & tlb_0_P0_V | tlbHit_1 & tlb_1_P0_V | tlbHit_2 & tlb_2_P0_V | tlbHit_3 & tlb_3_P0_V
     | tlbHit_4 & tlb_4_P0_V | tlbHit_5 & tlb_5_P0_V | tlbHit_6 & tlb_6_P0_V | tlbHit_7 & tlb_7_P0_V | tlbHit_8 &
    tlb_8_P0_V | tlbHit_9 & tlb_9_P0_V | tlbHit_10 & tlb_10_P0_V | tlbHit_11 & tlb_11_P0_V | tlbHit_12 & tlb_12_P0_V |
    tlbHit_13 & tlb_13_P0_V | tlbHit_14 & tlb_14_P0_V | _foundTLB_T_330;
  reg  tlb_16_P0_V;
  reg  tlb_17_P0_V;
  reg  tlb_18_P0_V;
  reg  tlb_19_P0_V;
  reg  tlb_20_P0_V;
  reg  tlb_21_P0_V;
  reg  tlb_22_P0_V;
  reg  tlb_23_P0_V;
  reg  tlb_24_P0_V;
  reg  tlb_25_P0_V;
  reg  tlb_26_P0_V;
  reg  tlb_27_P0_V;
  reg  tlb_28_P0_V;
  reg  tlb_29_P0_V;
  reg  tlb_30_P0_V;
  wire  _foundTLB_T_376 = _foundTLB_T_361 | tlbHit_16 & tlb_16_P0_V | tlbHit_17 & tlb_17_P0_V | tlbHit_18 & tlb_18_P0_V
     | tlbHit_19 & tlb_19_P0_V | tlbHit_20 & tlb_20_P0_V | tlbHit_21 & tlb_21_P0_V | tlbHit_22 & tlb_22_P0_V | tlbHit_23
     & tlb_23_P0_V | tlbHit_24 & tlb_24_P0_V | tlbHit_25 & tlb_25_P0_V | tlbHit_26 & tlb_26_P0_V | tlbHit_27 &
    tlb_27_P0_V | tlbHit_28 & tlb_28_P0_V | tlbHit_29 & tlb_29_P0_V | tlbHit_30 & tlb_30_P0_V;
  reg  tlb_31_P0_V;
  wire  foundTLB_P0_V = _foundTLB_T_376 | tlbHit_31 & tlb_31_P0_V;
  wire  foundP_V = oddPG ? foundTLB_P1_V : foundTLB_P0_V;
  wire  _GEN_11 = PC[31:29] == csrs_28_VSEG & (csrs_28_PLV0 & _T_11 | csrs_28_PLV3 & _T_13) ? 1'h0 : ~foundP_V;
  wire  invalid = PC[31:29] == csrs_27_VSEG & (csrs_27_PLV0 & crmd_PLV == 2'h0 | csrs_27_PLV3 & crmd_PLV == 2'h3) ? 1'h0
     : _GEN_11;
  reg [1:0] tlb_0_P1_PLV;
  wire [1:0] _foundTLB_T_189 = tlbHit_0 ? tlb_0_P1_PLV : 2'h0;
  reg [1:0] tlb_1_P1_PLV;
  wire [1:0] _foundTLB_T_190 = tlbHit_1 ? tlb_1_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_221 = _foundTLB_T_189 | _foundTLB_T_190;
  reg [1:0] tlb_2_P1_PLV;
  wire [1:0] _foundTLB_T_191 = tlbHit_2 ? tlb_2_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_222 = _foundTLB_T_221 | _foundTLB_T_191;
  reg [1:0] tlb_3_P1_PLV;
  wire [1:0] _foundTLB_T_192 = tlbHit_3 ? tlb_3_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_223 = _foundTLB_T_222 | _foundTLB_T_192;
  reg [1:0] tlb_4_P1_PLV;
  wire [1:0] _foundTLB_T_193 = tlbHit_4 ? tlb_4_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_224 = _foundTLB_T_223 | _foundTLB_T_193;
  reg [1:0] tlb_5_P1_PLV;
  wire [1:0] _foundTLB_T_194 = tlbHit_5 ? tlb_5_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_225 = _foundTLB_T_224 | _foundTLB_T_194;
  reg [1:0] tlb_6_P1_PLV;
  wire [1:0] _foundTLB_T_195 = tlbHit_6 ? tlb_6_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_226 = _foundTLB_T_225 | _foundTLB_T_195;
  reg [1:0] tlb_7_P1_PLV;
  wire [1:0] _foundTLB_T_196 = tlbHit_7 ? tlb_7_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_227 = _foundTLB_T_226 | _foundTLB_T_196;
  reg [1:0] tlb_8_P1_PLV;
  wire [1:0] _foundTLB_T_197 = tlbHit_8 ? tlb_8_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_228 = _foundTLB_T_227 | _foundTLB_T_197;
  reg [1:0] tlb_9_P1_PLV;
  wire [1:0] _foundTLB_T_198 = tlbHit_9 ? tlb_9_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_229 = _foundTLB_T_228 | _foundTLB_T_198;
  reg [1:0] tlb_10_P1_PLV;
  wire [1:0] _foundTLB_T_199 = tlbHit_10 ? tlb_10_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_230 = _foundTLB_T_229 | _foundTLB_T_199;
  reg [1:0] tlb_11_P1_PLV;
  wire [1:0] _foundTLB_T_200 = tlbHit_11 ? tlb_11_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_231 = _foundTLB_T_230 | _foundTLB_T_200;
  reg [1:0] tlb_12_P1_PLV;
  wire [1:0] _foundTLB_T_201 = tlbHit_12 ? tlb_12_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_232 = _foundTLB_T_231 | _foundTLB_T_201;
  reg [1:0] tlb_13_P1_PLV;
  wire [1:0] _foundTLB_T_202 = tlbHit_13 ? tlb_13_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_233 = _foundTLB_T_232 | _foundTLB_T_202;
  reg [1:0] tlb_14_P1_PLV;
  wire [1:0] _foundTLB_T_203 = tlbHit_14 ? tlb_14_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_234 = _foundTLB_T_233 | _foundTLB_T_203;
  reg [1:0] tlb_15_P1_PLV;
  wire [1:0] _foundTLB_T_204 = tlbHit_15 ? tlb_15_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_235 = _foundTLB_T_234 | _foundTLB_T_204;
  reg [1:0] tlb_16_P1_PLV;
  wire [1:0] _foundTLB_T_205 = tlbHit_16 ? tlb_16_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_236 = _foundTLB_T_235 | _foundTLB_T_205;
  reg [1:0] tlb_17_P1_PLV;
  wire [1:0] _foundTLB_T_206 = tlbHit_17 ? tlb_17_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_237 = _foundTLB_T_236 | _foundTLB_T_206;
  reg [1:0] tlb_18_P1_PLV;
  wire [1:0] _foundTLB_T_207 = tlbHit_18 ? tlb_18_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_238 = _foundTLB_T_237 | _foundTLB_T_207;
  reg [1:0] tlb_19_P1_PLV;
  wire [1:0] _foundTLB_T_208 = tlbHit_19 ? tlb_19_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_239 = _foundTLB_T_238 | _foundTLB_T_208;
  reg [1:0] tlb_20_P1_PLV;
  wire [1:0] _foundTLB_T_209 = tlbHit_20 ? tlb_20_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_240 = _foundTLB_T_239 | _foundTLB_T_209;
  reg [1:0] tlb_21_P1_PLV;
  wire [1:0] _foundTLB_T_210 = tlbHit_21 ? tlb_21_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_241 = _foundTLB_T_240 | _foundTLB_T_210;
  reg [1:0] tlb_22_P1_PLV;
  wire [1:0] _foundTLB_T_211 = tlbHit_22 ? tlb_22_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_242 = _foundTLB_T_241 | _foundTLB_T_211;
  reg [1:0] tlb_23_P1_PLV;
  wire [1:0] _foundTLB_T_212 = tlbHit_23 ? tlb_23_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_243 = _foundTLB_T_242 | _foundTLB_T_212;
  reg [1:0] tlb_24_P1_PLV;
  wire [1:0] _foundTLB_T_213 = tlbHit_24 ? tlb_24_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_244 = _foundTLB_T_243 | _foundTLB_T_213;
  reg [1:0] tlb_25_P1_PLV;
  wire [1:0] _foundTLB_T_214 = tlbHit_25 ? tlb_25_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_245 = _foundTLB_T_244 | _foundTLB_T_214;
  reg [1:0] tlb_26_P1_PLV;
  wire [1:0] _foundTLB_T_215 = tlbHit_26 ? tlb_26_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_246 = _foundTLB_T_245 | _foundTLB_T_215;
  reg [1:0] tlb_27_P1_PLV;
  wire [1:0] _foundTLB_T_216 = tlbHit_27 ? tlb_27_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_247 = _foundTLB_T_246 | _foundTLB_T_216;
  reg [1:0] tlb_28_P1_PLV;
  wire [1:0] _foundTLB_T_217 = tlbHit_28 ? tlb_28_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_248 = _foundTLB_T_247 | _foundTLB_T_217;
  reg [1:0] tlb_29_P1_PLV;
  wire [1:0] _foundTLB_T_218 = tlbHit_29 ? tlb_29_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_249 = _foundTLB_T_248 | _foundTLB_T_218;
  reg [1:0] tlb_30_P1_PLV;
  wire [1:0] _foundTLB_T_219 = tlbHit_30 ? tlb_30_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_250 = _foundTLB_T_249 | _foundTLB_T_219;
  reg [1:0] tlb_31_P1_PLV;
  wire [1:0] _foundTLB_T_220 = tlbHit_31 ? tlb_31_P1_PLV : 2'h0;
  wire [1:0] foundTLB_P1_PLV = _foundTLB_T_250 | _foundTLB_T_220;
  reg [1:0] tlb_0_P0_PLV;
  wire [1:0] _foundTLB_T_504 = tlbHit_0 ? tlb_0_P0_PLV : 2'h0;
  reg [1:0] tlb_1_P0_PLV;
  wire [1:0] _foundTLB_T_505 = tlbHit_1 ? tlb_1_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_536 = _foundTLB_T_504 | _foundTLB_T_505;
  reg [1:0] tlb_2_P0_PLV;
  wire [1:0] _foundTLB_T_506 = tlbHit_2 ? tlb_2_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_537 = _foundTLB_T_536 | _foundTLB_T_506;
  reg [1:0] tlb_3_P0_PLV;
  wire [1:0] _foundTLB_T_507 = tlbHit_3 ? tlb_3_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_538 = _foundTLB_T_537 | _foundTLB_T_507;
  reg [1:0] tlb_4_P0_PLV;
  wire [1:0] _foundTLB_T_508 = tlbHit_4 ? tlb_4_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_539 = _foundTLB_T_538 | _foundTLB_T_508;
  reg [1:0] tlb_5_P0_PLV;
  wire [1:0] _foundTLB_T_509 = tlbHit_5 ? tlb_5_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_540 = _foundTLB_T_539 | _foundTLB_T_509;
  reg [1:0] tlb_6_P0_PLV;
  wire [1:0] _foundTLB_T_510 = tlbHit_6 ? tlb_6_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_541 = _foundTLB_T_540 | _foundTLB_T_510;
  reg [1:0] tlb_7_P0_PLV;
  wire [1:0] _foundTLB_T_511 = tlbHit_7 ? tlb_7_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_542 = _foundTLB_T_541 | _foundTLB_T_511;
  reg [1:0] tlb_8_P0_PLV;
  wire [1:0] _foundTLB_T_512 = tlbHit_8 ? tlb_8_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_543 = _foundTLB_T_542 | _foundTLB_T_512;
  reg [1:0] tlb_9_P0_PLV;
  wire [1:0] _foundTLB_T_513 = tlbHit_9 ? tlb_9_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_544 = _foundTLB_T_543 | _foundTLB_T_513;
  reg [1:0] tlb_10_P0_PLV;
  wire [1:0] _foundTLB_T_514 = tlbHit_10 ? tlb_10_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_545 = _foundTLB_T_544 | _foundTLB_T_514;
  reg [1:0] tlb_11_P0_PLV;
  wire [1:0] _foundTLB_T_515 = tlbHit_11 ? tlb_11_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_546 = _foundTLB_T_545 | _foundTLB_T_515;
  reg [1:0] tlb_12_P0_PLV;
  wire [1:0] _foundTLB_T_516 = tlbHit_12 ? tlb_12_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_547 = _foundTLB_T_546 | _foundTLB_T_516;
  reg [1:0] tlb_13_P0_PLV;
  wire [1:0] _foundTLB_T_517 = tlbHit_13 ? tlb_13_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_548 = _foundTLB_T_547 | _foundTLB_T_517;
  reg [1:0] tlb_14_P0_PLV;
  wire [1:0] _foundTLB_T_518 = tlbHit_14 ? tlb_14_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_549 = _foundTLB_T_548 | _foundTLB_T_518;
  reg [1:0] tlb_15_P0_PLV;
  wire [1:0] _foundTLB_T_519 = tlbHit_15 ? tlb_15_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_550 = _foundTLB_T_549 | _foundTLB_T_519;
  reg [1:0] tlb_16_P0_PLV;
  wire [1:0] _foundTLB_T_520 = tlbHit_16 ? tlb_16_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_551 = _foundTLB_T_550 | _foundTLB_T_520;
  reg [1:0] tlb_17_P0_PLV;
  wire [1:0] _foundTLB_T_521 = tlbHit_17 ? tlb_17_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_552 = _foundTLB_T_551 | _foundTLB_T_521;
  reg [1:0] tlb_18_P0_PLV;
  wire [1:0] _foundTLB_T_522 = tlbHit_18 ? tlb_18_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_553 = _foundTLB_T_552 | _foundTLB_T_522;
  reg [1:0] tlb_19_P0_PLV;
  wire [1:0] _foundTLB_T_523 = tlbHit_19 ? tlb_19_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_554 = _foundTLB_T_553 | _foundTLB_T_523;
  reg [1:0] tlb_20_P0_PLV;
  wire [1:0] _foundTLB_T_524 = tlbHit_20 ? tlb_20_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_555 = _foundTLB_T_554 | _foundTLB_T_524;
  reg [1:0] tlb_21_P0_PLV;
  wire [1:0] _foundTLB_T_525 = tlbHit_21 ? tlb_21_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_556 = _foundTLB_T_555 | _foundTLB_T_525;
  reg [1:0] tlb_22_P0_PLV;
  wire [1:0] _foundTLB_T_526 = tlbHit_22 ? tlb_22_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_557 = _foundTLB_T_556 | _foundTLB_T_526;
  reg [1:0] tlb_23_P0_PLV;
  wire [1:0] _foundTLB_T_527 = tlbHit_23 ? tlb_23_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_558 = _foundTLB_T_557 | _foundTLB_T_527;
  reg [1:0] tlb_24_P0_PLV;
  wire [1:0] _foundTLB_T_528 = tlbHit_24 ? tlb_24_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_559 = _foundTLB_T_558 | _foundTLB_T_528;
  reg [1:0] tlb_25_P0_PLV;
  wire [1:0] _foundTLB_T_529 = tlbHit_25 ? tlb_25_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_560 = _foundTLB_T_559 | _foundTLB_T_529;
  reg [1:0] tlb_26_P0_PLV;
  wire [1:0] _foundTLB_T_530 = tlbHit_26 ? tlb_26_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_561 = _foundTLB_T_560 | _foundTLB_T_530;
  reg [1:0] tlb_27_P0_PLV;
  wire [1:0] _foundTLB_T_531 = tlbHit_27 ? tlb_27_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_562 = _foundTLB_T_561 | _foundTLB_T_531;
  reg [1:0] tlb_28_P0_PLV;
  wire [1:0] _foundTLB_T_532 = tlbHit_28 ? tlb_28_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_563 = _foundTLB_T_562 | _foundTLB_T_532;
  reg [1:0] tlb_29_P0_PLV;
  wire [1:0] _foundTLB_T_533 = tlbHit_29 ? tlb_29_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_564 = _foundTLB_T_563 | _foundTLB_T_533;
  reg [1:0] tlb_30_P0_PLV;
  wire [1:0] _foundTLB_T_534 = tlbHit_30 ? tlb_30_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_565 = _foundTLB_T_564 | _foundTLB_T_534;
  reg [1:0] tlb_31_P0_PLV;
  wire [1:0] _foundTLB_T_535 = tlbHit_31 ? tlb_31_P0_PLV : 2'h0;
  wire [1:0] foundTLB_P0_PLV = _foundTLB_T_565 | _foundTLB_T_535;
  wire [1:0] foundP_PLV = oddPG ? foundTLB_P1_PLV : foundTLB_P0_PLV;
  wire  _GEN_12 = PC[31:29] == csrs_28_VSEG & (csrs_28_PLV0 & _T_11 | csrs_28_PLV3 & _T_13) ? 1'h0 : crmd_PLV >
    foundP_PLV;
  wire  ppi = PC[31:29] == csrs_27_VSEG & (csrs_27_PLV0 & crmd_PLV == 2'h0 | csrs_27_PLV3 & crmd_PLV == 2'h3) ? 1'h0 :
    _GEN_12;
  wire  _GEN_21 = ppi ? 1'h0 : 1'h1;
  wire  _GEN_24 = invalid ? 1'h0 : _GEN_21;
  wire  _GEN_28 = miss ? 1'h0 : _GEN_24;
  wire  _GEN_29 = crmd_DA | _GEN_28;
  wire  _GEN_34 = PC[1:0] != 2'h0 | PC[31] & crmd_PLV != 2'h0 ? 1'h0 : _GEN_29;
  wire  _GEN_39 = ~INT & ~idle & _GEN_34;
  wire  IF_OK = dStallReg | iStallReg | _GEN_39;
  wire  iStall = ~io_inst_resp_valid & (io_inst_req_valid | iStallReg);
  wire  _T_1319 = ~iStall;
  reg [31:0] inst_reg;
  wire [31:0] inst = dStallReg ? inst_reg : io_inst_resp_bits;
  wire [31:0] _T_37 = inst & 32'hfffffc1f;
  wire  _T_38 = 32'h6000 == _T_37;
  wire [31:0] _T_39 = inst & 32'hffffffe0;
  wire  _T_40 = 32'h6000 == _T_39;
  wire  _T_42 = 32'h6400 == _T_39;
  wire [31:0] _T_43 = inst & 32'hffff8000;
  wire  _T_44 = 32'h100000 == _T_43;
  wire  _T_46 = 32'h110000 == _T_43;
  wire  _T_48 = 32'h120000 == _T_43;
  wire  _T_50 = 32'h128000 == _T_43;
  wire  _T_52 = 32'h140000 == _T_43;
  wire  _T_54 = 32'h148000 == _T_43;
  wire  _T_56 = 32'h150000 == _T_43;
  wire  _T_58 = 32'h158000 == _T_43;
  wire  _T_60 = 32'h170000 == _T_43;
  wire  _T_62 = 32'h178000 == _T_43;
  wire  _T_64 = 32'h180000 == _T_43;
  wire  _T_66 = 32'h1c0000 == _T_43;
  wire  _T_68 = 32'h1c8000 == _T_43;
  wire  _T_70 = 32'h1d0000 == _T_43;
  wire  _T_72 = 32'h200000 == _T_43;
  wire  _T_74 = 32'h208000 == _T_43;
  wire  _T_76 = 32'h210000 == _T_43;
  wire  _T_78 = 32'h218000 == _T_43;
  wire  _T_80 = 32'h2a0000 == _T_43;
  wire  _T_82 = 32'h2b0000 == _T_43;
  wire  _T_84 = 32'h408000 == _T_43;
  wire  _T_86 = 32'h448000 == _T_43;
  wire  _T_88 = 32'h488000 == _T_43;
  wire [31:0] _T_89 = inst & 32'hffc00000;
  wire  _T_90 = 32'h2000000 == _T_89;
  wire  _T_92 = 32'h2400000 == _T_89;
  wire  _T_94 = 32'h2800000 == _T_89;
  wire  _T_96 = 32'h3400000 == _T_89;
  wire  _T_98 = 32'h3800000 == _T_89;
  wire  _T_100 = 32'h3c00000 == _T_89;
  wire [31:0] _T_101 = inst & 32'hff000000;
  wire  _T_102 = 32'h4000000 == _T_101;
  wire  _T_104 = 32'h6000000 == _T_89;
  wire  _T_106 = 32'h6482800 == inst;
  wire  _T_108 = 32'h6482c00 == inst;
  wire  _T_110 = 32'h6483000 == inst;
  wire  _T_112 = 32'h6483400 == inst;
  wire  _T_114 = 32'h6498000 == _T_43;
  wire  _T_116 = 32'h6483800 == inst;
  wire  _T_118 = 32'h6488000 == _T_43;
  wire [31:0] _T_119 = inst & 32'hfe000000;
  wire  _T_120 = 32'h14000000 == _T_119;
  wire  _T_122 = 32'h1c000000 == _T_119;
  wire  _T_124 = 32'h20000000 == _T_101;
  wire  _T_126 = 32'h21000000 == _T_101;
  wire  _T_128 = 32'h28000000 == _T_89;
  wire  _T_130 = 32'h28400000 == _T_89;
  wire  _T_132 = 32'h28800000 == _T_89;
  wire  _T_134 = 32'h29000000 == _T_89;
  wire  _T_136 = 32'h29400000 == _T_89;
  wire  _T_138 = 32'h29800000 == _T_89;
  wire  _T_140 = 32'h2a000000 == _T_89;
  wire  _T_142 = 32'h2a400000 == _T_89;
  wire  _T_144 = 32'h2ac00000 == _T_89;
  wire  _T_146 = 32'h38720000 == _T_43;
  wire  _T_148 = 32'h38728000 == _T_43;
  wire [31:0] _T_149 = inst & 32'hfc000000;
  wire  _T_150 = 32'h4c000000 == _T_149;
  wire  _T_152 = 32'h50000000 == _T_149;
  wire  _T_154 = 32'h54000000 == _T_149;
  wire  _T_156 = 32'h58000000 == _T_149;
  wire  _T_158 = 32'h5c000000 == _T_149;
  wire  _T_160 = 32'h60000000 == _T_149;
  wire  _T_162 = 32'h64000000 == _T_149;
  wire  _T_164 = 32'h68000000 == _T_149;
  wire  _T_166 = 32'h6c000000 == _T_149;
  wire  _T_914 = _T_80 ? 1'h0 : _T_82;
  wire  _T_915 = _T_78 ? 1'h0 : _T_914;
  wire  _T_916 = _T_76 ? 1'h0 : _T_915;
  wire  _T_917 = _T_74 ? 1'h0 : _T_916;
  wire  _T_918 = _T_72 ? 1'h0 : _T_917;
  wire  _T_919 = _T_70 ? 1'h0 : _T_918;
  wire  _T_920 = _T_68 ? 1'h0 : _T_919;
  wire  _T_921 = _T_66 ? 1'h0 : _T_920;
  wire  _T_922 = _T_64 ? 1'h0 : _T_921;
  wire  _T_923 = _T_62 ? 1'h0 : _T_922;
  wire  _T_924 = _T_60 ? 1'h0 : _T_923;
  wire  _T_925 = _T_58 ? 1'h0 : _T_924;
  wire  _T_926 = _T_56 ? 1'h0 : _T_925;
  wire  _T_927 = _T_54 ? 1'h0 : _T_926;
  wire  _T_928 = _T_52 ? 1'h0 : _T_927;
  wire  _T_929 = _T_50 ? 1'h0 : _T_928;
  wire  _T_930 = _T_48 ? 1'h0 : _T_929;
  wire  _T_931 = _T_46 ? 1'h0 : _T_930;
  wire  _T_932 = _T_44 ? 1'h0 : _T_931;
  wire  _T_933 = _T_42 ? 1'h0 : _T_932;
  wire  _T_934 = _T_40 ? 1'h0 : _T_933;
  wire  c0_6 = _T_38 ? 1'h0 : _T_934;
  wire  _T_851 = _T_78 ? 1'h0 : _T_80;
  wire  _T_852 = _T_76 ? 1'h0 : _T_851;
  wire  _T_853 = _T_74 ? 1'h0 : _T_852;
  wire  _T_854 = _T_72 ? 1'h0 : _T_853;
  wire  _T_855 = _T_70 ? 1'h0 : _T_854;
  wire  _T_856 = _T_68 ? 1'h0 : _T_855;
  wire  _T_857 = _T_66 ? 1'h0 : _T_856;
  wire  _T_858 = _T_64 ? 1'h0 : _T_857;
  wire  _T_859 = _T_62 ? 1'h0 : _T_858;
  wire  _T_860 = _T_60 ? 1'h0 : _T_859;
  wire  _T_861 = _T_58 ? 1'h0 : _T_860;
  wire  _T_862 = _T_56 ? 1'h0 : _T_861;
  wire  _T_863 = _T_54 ? 1'h0 : _T_862;
  wire  _T_864 = _T_52 ? 1'h0 : _T_863;
  wire  _T_865 = _T_50 ? 1'h0 : _T_864;
  wire  _T_866 = _T_48 ? 1'h0 : _T_865;
  wire  _T_867 = _T_46 ? 1'h0 : _T_866;
  wire  _T_868 = _T_44 ? 1'h0 : _T_867;
  wire  _T_869 = _T_42 ? 1'h0 : _T_868;
  wire  _T_870 = _T_40 ? 1'h0 : _T_869;
  wire  break_ = _T_38 ? 1'h0 : _T_870;
  wire  _T_197 = _T_106 | (_T_108 | (_T_110 | (_T_112 | (_T_114 | (_T_116 | (_T_118 | (_T_120 | (_T_122 | (_T_124 | (
    _T_126 | (_T_128 | (_T_130 | (_T_132 | (_T_134 | (_T_136 | (_T_138 | (_T_140 | (_T_142 | (_T_144 | (_T_146 | (_T_148
     | (_T_150 | (_T_152 | (_T_154 | (_T_156 | (_T_158 | (_T_160 | (_T_162 | (_T_164 | _T_166)))))))))))))))))))))))))))
    ));
  wire  _T_227 = _T_46 | (_T_48 | (_T_50 | (_T_52 | (_T_54 | (_T_56 | (_T_58 | (_T_60 | (_T_62 | (_T_64 | (_T_66 | (
    _T_68 | (_T_70 | (_T_72 | (_T_74 | (_T_76 | (_T_78 | (_T_80 | (_T_82 | (_T_84 | (_T_86 | (_T_88 | (_T_90 | (_T_92 |
    (_T_94 | (_T_96 | (_T_98 | (_T_100 | (_T_102 | (_T_104 | _T_197)))))))))))))))))))))))))))));
  wire  instV = _T_38 | (_T_40 | (_T_42 | (_T_44 | _T_227)));
  wire  _T_1324 = ~c0_6 & ~break_ & instV;
  wire  _GEN_55 = IF_OK & ~iStall & _T_1324;
  wire  ID_OK = dStallReg | _GEN_55;
  wire [2:0] _T_690 = _T_144 ? 3'h0 : 3'h7;
  wire [2:0] _T_691 = _T_142 ? 3'h3 : _T_690;
  wire [2:0] _T_692 = _T_140 ? 3'h1 : _T_691;
  wire [2:0] _T_693 = _T_138 ? 3'h4 : _T_692;
  wire [2:0] _T_694 = _T_136 ? 3'h2 : _T_693;
  wire [2:0] _T_695 = _T_134 ? 3'h0 : _T_694;
  wire [2:0] _T_696 = _T_132 ? 3'h4 : _T_695;
  wire [2:0] _T_697 = _T_130 ? 3'h2 : _T_696;
  wire [2:0] _T_698 = _T_128 ? 3'h0 : _T_697;
  wire [2:0] _T_699 = _T_126 ? 3'h4 : _T_698;
  wire [2:0] _T_700 = _T_124 ? 3'h4 : _T_699;
  wire [2:0] _T_701 = _T_122 ? 3'h7 : _T_700;
  wire [2:0] _T_702 = _T_120 ? 3'h7 : _T_701;
  wire [2:0] _T_703 = _T_118 ? 3'h7 : _T_702;
  wire [2:0] _T_704 = _T_116 ? 3'h7 : _T_703;
  wire [2:0] _T_705 = _T_114 ? 3'h7 : _T_704;
  wire [2:0] _T_706 = _T_112 ? 3'h7 : _T_705;
  wire [2:0] _T_707 = _T_110 ? 3'h7 : _T_706;
  wire [2:0] _T_708 = _T_108 ? 3'h7 : _T_707;
  wire [2:0] _T_709 = _T_106 ? 3'h7 : _T_708;
  wire [2:0] _T_710 = _T_104 ? 3'h0 : _T_709;
  wire [2:0] _T_711 = _T_102 ? 3'h7 : _T_710;
  wire [2:0] _T_712 = _T_100 ? 3'h7 : _T_711;
  wire [2:0] _T_713 = _T_98 ? 3'h7 : _T_712;
  wire [2:0] _T_714 = _T_96 ? 3'h7 : _T_713;
  wire [2:0] _T_715 = _T_94 ? 3'h7 : _T_714;
  wire [2:0] _T_716 = _T_92 ? 3'h7 : _T_715;
  wire [2:0] _T_717 = _T_90 ? 3'h7 : _T_716;
  wire [2:0] _T_718 = _T_88 ? 3'h7 : _T_717;
  wire [2:0] _T_719 = _T_86 ? 3'h7 : _T_718;
  wire [2:0] _T_720 = _T_84 ? 3'h7 : _T_719;
  wire [2:0] _T_721 = _T_82 ? 3'h7 : _T_720;
  wire [2:0] _T_722 = _T_80 ? 3'h7 : _T_721;
  wire [2:0] _T_723 = _T_78 ? 3'h7 : _T_722;
  wire [2:0] _T_724 = _T_76 ? 3'h7 : _T_723;
  wire [2:0] _T_725 = _T_74 ? 3'h7 : _T_724;
  wire [2:0] _T_726 = _T_72 ? 3'h7 : _T_725;
  wire [2:0] _T_727 = _T_70 ? 3'h7 : _T_726;
  wire [2:0] _T_728 = _T_68 ? 3'h7 : _T_727;
  wire [2:0] _T_729 = _T_66 ? 3'h7 : _T_728;
  wire [2:0] _T_730 = _T_64 ? 3'h7 : _T_729;
  wire [2:0] _T_731 = _T_62 ? 3'h7 : _T_730;
  wire [2:0] _T_732 = _T_60 ? 3'h7 : _T_731;
  wire [2:0] _T_733 = _T_58 ? 3'h7 : _T_732;
  wire [2:0] _T_734 = _T_56 ? 3'h7 : _T_733;
  wire [2:0] _T_735 = _T_54 ? 3'h7 : _T_734;
  wire [2:0] _T_736 = _T_52 ? 3'h7 : _T_735;
  wire [2:0] _T_737 = _T_50 ? 3'h7 : _T_736;
  wire [2:0] _T_738 = _T_48 ? 3'h7 : _T_737;
  wire [2:0] _T_739 = _T_46 ? 3'h7 : _T_738;
  wire [2:0] _T_740 = _T_44 ? 3'h7 : _T_739;
  wire [2:0] _T_741 = _T_42 ? 3'h7 : _T_740;
  wire [2:0] _T_742 = _T_40 ? 3'h7 : _T_741;
  wire [2:0] c0_3 = _T_38 ? 3'h7 : _T_742;
  wire  _T_1223 = _T_102 ? 1'h0 : _T_104;
  wire  _T_1224 = _T_100 ? 1'h0 : _T_1223;
  wire  _T_1225 = _T_98 ? 1'h0 : _T_1224;
  wire  _T_1226 = _T_96 ? 1'h0 : _T_1225;
  wire  _T_1227 = _T_94 ? 1'h0 : _T_1226;
  wire  _T_1228 = _T_92 ? 1'h0 : _T_1227;
  wire  _T_1229 = _T_90 ? 1'h0 : _T_1228;
  wire  _T_1230 = _T_88 ? 1'h0 : _T_1229;
  wire  _T_1231 = _T_86 ? 1'h0 : _T_1230;
  wire  _T_1232 = _T_84 ? 1'h0 : _T_1231;
  wire  _T_1233 = _T_82 ? 1'h0 : _T_1232;
  wire  _T_1234 = _T_80 ? 1'h0 : _T_1233;
  wire  _T_1235 = _T_78 ? 1'h0 : _T_1234;
  wire  _T_1236 = _T_76 ? 1'h0 : _T_1235;
  wire  _T_1237 = _T_74 ? 1'h0 : _T_1236;
  wire  _T_1238 = _T_72 ? 1'h0 : _T_1237;
  wire  _T_1239 = _T_70 ? 1'h0 : _T_1238;
  wire  _T_1240 = _T_68 ? 1'h0 : _T_1239;
  wire  _T_1241 = _T_66 ? 1'h0 : _T_1240;
  wire  _T_1242 = _T_64 ? 1'h0 : _T_1241;
  wire  _T_1243 = _T_62 ? 1'h0 : _T_1242;
  wire  _T_1244 = _T_60 ? 1'h0 : _T_1243;
  wire  _T_1245 = _T_58 ? 1'h0 : _T_1244;
  wire  _T_1246 = _T_56 ? 1'h0 : _T_1245;
  wire  _T_1247 = _T_54 ? 1'h0 : _T_1246;
  wire  _T_1248 = _T_52 ? 1'h0 : _T_1247;
  wire  _T_1249 = _T_50 ? 1'h0 : _T_1248;
  wire  _T_1250 = _T_48 ? 1'h0 : _T_1249;
  wire  _T_1251 = _T_46 ? 1'h0 : _T_1250;
  wire  _T_1252 = _T_44 ? 1'h0 : _T_1251;
  wire  _T_1253 = _T_42 ? 1'h0 : _T_1252;
  wire  _T_1254 = _T_40 ? 1'h0 : _T_1253;
  wire  c0_11 = _T_38 ? 1'h0 : _T_1254;
  wire [4:0] d = inst[4:0];
  wire [4:0] _T_423 = _T_166 ? 5'h0 : 5'h13;
  wire [4:0] _T_424 = _T_164 ? 5'h0 : _T_423;
  wire [4:0] _T_425 = _T_162 ? 5'h0 : _T_424;
  wire [4:0] _T_426 = _T_160 ? 5'h0 : _T_425;
  wire [4:0] _T_427 = _T_158 ? 5'h0 : _T_426;
  wire [4:0] _T_428 = _T_156 ? 5'h0 : _T_427;
  wire [4:0] _T_429 = _T_154 ? 5'h0 : _T_428;
  wire [4:0] _T_430 = _T_152 ? 5'h0 : _T_429;
  wire [4:0] _T_431 = _T_150 ? 5'h0 : _T_430;
  wire [4:0] _T_432 = _T_148 ? 5'h13 : _T_431;
  wire [4:0] _T_433 = _T_146 ? 5'h13 : _T_432;
  wire [4:0] _T_434 = _T_144 ? 5'h0 : _T_433;
  wire [4:0] _T_435 = _T_142 ? 5'h0 : _T_434;
  wire [4:0] _T_436 = _T_140 ? 5'h0 : _T_435;
  wire [4:0] _T_437 = _T_138 ? 5'h0 : _T_436;
  wire [4:0] _T_438 = _T_136 ? 5'h0 : _T_437;
  wire [4:0] _T_439 = _T_134 ? 5'h0 : _T_438;
  wire [4:0] _T_440 = _T_132 ? 5'h0 : _T_439;
  wire [4:0] _T_441 = _T_130 ? 5'h0 : _T_440;
  wire [4:0] _T_442 = _T_128 ? 5'h0 : _T_441;
  wire [4:0] _T_443 = _T_126 ? 5'h0 : _T_442;
  wire [4:0] _T_444 = _T_124 ? 5'h0 : _T_443;
  wire [4:0] _T_445 = _T_122 ? 5'h0 : _T_444;
  wire [4:0] _T_446 = _T_120 ? 5'hb : _T_445;
  wire [4:0] _T_447 = _T_118 ? 5'h13 : _T_446;
  wire [4:0] _T_448 = _T_116 ? 5'h13 : _T_447;
  wire [4:0] _T_449 = _T_114 ? 5'h13 : _T_448;
  wire [4:0] _T_450 = _T_112 ? 5'h13 : _T_449;
  wire [4:0] _T_451 = _T_110 ? 5'h13 : _T_450;
  wire [4:0] _T_452 = _T_108 ? 5'h13 : _T_451;
  wire [4:0] _T_453 = _T_106 ? 5'h13 : _T_452;
  wire [4:0] _T_454 = _T_104 ? 5'h0 : _T_453;
  wire [4:0] _T_455 = _T_102 ? 5'h13 : _T_454;
  wire [4:0] _T_456 = _T_100 ? 5'h8 : _T_455;
  wire [4:0] _T_457 = _T_98 ? 5'h6 : _T_456;
  wire [4:0] _T_458 = _T_96 ? 5'h5 : _T_457;
  wire [4:0] _T_459 = _T_94 ? 5'h0 : _T_458;
  wire [4:0] _T_460 = _T_92 ? 5'ha : _T_459;
  wire [4:0] _T_461 = _T_90 ? 5'h9 : _T_460;
  wire [4:0] _T_462 = _T_88 ? 5'h4 : _T_461;
  wire [4:0] _T_463 = _T_86 ? 5'h3 : _T_462;
  wire [4:0] _T_464 = _T_84 ? 5'h2 : _T_463;
  wire [4:0] _T_465 = _T_82 ? 5'h13 : _T_464;
  wire [4:0] _T_466 = _T_80 ? 5'h13 : _T_465;
  wire [4:0] _T_467 = _T_78 ? 5'h11 : _T_466;
  wire [4:0] _T_468 = _T_76 ? 5'h12 : _T_467;
  wire [4:0] _T_469 = _T_74 ? 5'hf : _T_468;
  wire [4:0] _T_470 = _T_72 ? 5'h10 : _T_469;
  wire [4:0] _T_471 = _T_70 ? 5'he : _T_470;
  wire [4:0] _T_472 = _T_68 ? 5'hd : _T_471;
  wire [4:0] _T_473 = _T_66 ? 5'hc : _T_472;
  wire [4:0] _T_474 = _T_64 ? 5'h4 : _T_473;
  wire [4:0] _T_475 = _T_62 ? 5'h3 : _T_474;
  wire [4:0] _T_476 = _T_60 ? 5'h2 : _T_475;
  wire [4:0] _T_477 = _T_58 ? 5'h8 : _T_476;
  wire [4:0] _T_478 = _T_56 ? 5'h6 : _T_477;
  wire [4:0] _T_479 = _T_54 ? 5'h5 : _T_478;
  wire [4:0] _T_480 = _T_52 ? 5'h7 : _T_479;
  wire [4:0] _T_481 = _T_50 ? 5'ha : _T_480;
  wire [4:0] _T_482 = _T_48 ? 5'h9 : _T_481;
  wire [4:0] _T_483 = _T_46 ? 5'h1 : _T_482;
  wire [4:0] _T_484 = _T_44 ? 5'h0 : _T_483;
  wire [4:0] _T_485 = _T_42 ? 5'h13 : _T_484;
  wire [4:0] _T_486 = _T_40 ? 5'h13 : _T_485;
  wire [4:0] func = _T_38 ? 5'h13 : _T_486;
  wire  _aluOut_T = func == 5'h0;
  wire  _T_303 = _T_150 ? 1'h0 : _T_152 | (_T_154 | (_T_156 | (_T_158 | (_T_160 | (_T_162 | (_T_164 | _T_166))))));
  wire  _T_304 = _T_148 ? 1'h0 : _T_303;
  wire  _T_305 = _T_146 ? 1'h0 : _T_304;
  wire  _T_306 = _T_144 ? 1'h0 : _T_305;
  wire  _T_307 = _T_142 ? 1'h0 : _T_306;
  wire  _T_308 = _T_140 ? 1'h0 : _T_307;
  wire  _T_309 = _T_138 ? 1'h0 : _T_308;
  wire  _T_310 = _T_136 ? 1'h0 : _T_309;
  wire  _T_311 = _T_134 ? 1'h0 : _T_310;
  wire  _T_312 = _T_132 ? 1'h0 : _T_311;
  wire  _T_313 = _T_130 ? 1'h0 : _T_312;
  wire  _T_314 = _T_128 ? 1'h0 : _T_313;
  wire  _T_315 = _T_126 ? 1'h0 : _T_314;
  wire  _T_316 = _T_124 ? 1'h0 : _T_315;
  wire  _T_318 = _T_120 ? 1'h0 : _T_122 | _T_316;
  wire  _T_319 = _T_118 ? 1'h0 : _T_318;
  wire  _T_320 = _T_116 ? 1'h0 : _T_319;
  wire  _T_321 = _T_114 ? 1'h0 : _T_320;
  wire  _T_322 = _T_112 ? 1'h0 : _T_321;
  wire  _T_323 = _T_110 ? 1'h0 : _T_322;
  wire  _T_324 = _T_108 ? 1'h0 : _T_323;
  wire  _T_325 = _T_106 ? 1'h0 : _T_324;
  wire  _T_326 = _T_104 ? 1'h0 : _T_325;
  wire  _T_327 = _T_102 ? 1'h0 : _T_326;
  wire  _T_328 = _T_100 ? 1'h0 : _T_327;
  wire  _T_329 = _T_98 ? 1'h0 : _T_328;
  wire  _T_330 = _T_96 ? 1'h0 : _T_329;
  wire  _T_331 = _T_94 ? 1'h0 : _T_330;
  wire  _T_332 = _T_92 ? 1'h0 : _T_331;
  wire  _T_333 = _T_90 ? 1'h0 : _T_332;
  wire  _T_334 = _T_88 ? 1'h0 : _T_333;
  wire  _T_335 = _T_86 ? 1'h0 : _T_334;
  wire  _T_336 = _T_84 ? 1'h0 : _T_335;
  wire  _T_337 = _T_82 ? 1'h0 : _T_336;
  wire  _T_338 = _T_80 ? 1'h0 : _T_337;
  wire  _T_339 = _T_78 ? 1'h0 : _T_338;
  wire  _T_340 = _T_76 ? 1'h0 : _T_339;
  wire  _T_341 = _T_74 ? 1'h0 : _T_340;
  wire  _T_342 = _T_72 ? 1'h0 : _T_341;
  wire  _T_343 = _T_70 ? 1'h0 : _T_342;
  wire  _T_344 = _T_68 ? 1'h0 : _T_343;
  wire  _T_345 = _T_66 ? 1'h0 : _T_344;
  wire  _T_346 = _T_64 ? 1'h0 : _T_345;
  wire  _T_347 = _T_62 ? 1'h0 : _T_346;
  wire  _T_348 = _T_60 ? 1'h0 : _T_347;
  wire  _T_349 = _T_58 ? 1'h0 : _T_348;
  wire  _T_350 = _T_56 ? 1'h0 : _T_349;
  wire  _T_351 = _T_54 ? 1'h0 : _T_350;
  wire  _T_352 = _T_52 ? 1'h0 : _T_351;
  wire  _T_353 = _T_50 ? 1'h0 : _T_352;
  wire  _T_354 = _T_48 ? 1'h0 : _T_353;
  wire  _T_355 = _T_46 ? 1'h0 : _T_354;
  wire  _T_356 = _T_44 ? 1'h0 : _T_355;
  wire  _T_357 = _T_42 ? 1'h0 : _T_356;
  wire  _T_358 = _T_40 ? 1'h0 : _T_357;
  wire  op1Sel = _T_38 ? 1'h0 : _T_358;
  wire [4:0] j = inst[9:5];
  wire [31:0] rj = j == 5'h0 ? 32'h0 : GR_rj_MPORT_data;
  wire [31:0] aluOp1 = ~op1Sel ? rj : PC;
  wire [2:0] _T_359 = _T_166 ? 3'h5 : 3'h0;
  wire [2:0] _T_360 = _T_164 ? 3'h5 : _T_359;
  wire [2:0] _T_361 = _T_162 ? 3'h5 : _T_360;
  wire [2:0] _T_362 = _T_160 ? 3'h5 : _T_361;
  wire [2:0] _T_363 = _T_158 ? 3'h5 : _T_362;
  wire [2:0] _T_364 = _T_156 ? 3'h5 : _T_363;
  wire [2:0] _T_365 = _T_154 ? 3'h7 : _T_364;
  wire [2:0] _T_366 = _T_152 ? 3'h7 : _T_365;
  wire [2:0] _T_367 = _T_150 ? 3'h5 : _T_366;
  wire [2:0] _T_368 = _T_148 ? 3'h0 : _T_367;
  wire [2:0] _T_369 = _T_146 ? 3'h0 : _T_368;
  wire [2:0] _T_370 = _T_144 ? 3'h3 : _T_369;
  wire [2:0] _T_371 = _T_142 ? 3'h3 : _T_370;
  wire [2:0] _T_372 = _T_140 ? 3'h3 : _T_371;
  wire [2:0] _T_373 = _T_138 ? 3'h3 : _T_372;
  wire [2:0] _T_374 = _T_136 ? 3'h3 : _T_373;
  wire [2:0] _T_375 = _T_134 ? 3'h3 : _T_374;
  wire [2:0] _T_376 = _T_132 ? 3'h3 : _T_375;
  wire [2:0] _T_377 = _T_130 ? 3'h3 : _T_376;
  wire [2:0] _T_378 = _T_128 ? 3'h3 : _T_377;
  wire [2:0] _T_379 = _T_126 ? 3'h4 : _T_378;
  wire [2:0] _T_380 = _T_124 ? 3'h4 : _T_379;
  wire [2:0] _T_381 = _T_122 ? 3'h6 : _T_380;
  wire [2:0] _T_382 = _T_120 ? 3'h6 : _T_381;
  wire [2:0] _T_383 = _T_118 ? 3'h0 : _T_382;
  wire [2:0] _T_384 = _T_116 ? 3'h0 : _T_383;
  wire [2:0] _T_385 = _T_114 ? 3'h0 : _T_384;
  wire [2:0] _T_386 = _T_112 ? 3'h0 : _T_385;
  wire [2:0] _T_387 = _T_110 ? 3'h0 : _T_386;
  wire [2:0] _T_388 = _T_108 ? 3'h0 : _T_387;
  wire [2:0] _T_389 = _T_106 ? 3'h0 : _T_388;
  wire [2:0] _T_390 = _T_104 ? 3'h3 : _T_389;
  wire [2:0] _T_391 = _T_102 ? 3'h0 : _T_390;
  wire [2:0] _T_392 = _T_100 ? 3'h2 : _T_391;
  wire [2:0] _T_393 = _T_98 ? 3'h2 : _T_392;
  wire [2:0] _T_394 = _T_96 ? 3'h2 : _T_393;
  wire [2:0] _T_395 = _T_94 ? 3'h3 : _T_394;
  wire [2:0] _T_396 = _T_92 ? 3'h3 : _T_395;
  wire [2:0] _T_397 = _T_90 ? 3'h3 : _T_396;
  wire [2:0] _T_398 = _T_88 ? 3'h1 : _T_397;
  wire [2:0] _T_399 = _T_86 ? 3'h1 : _T_398;
  wire [2:0] _T_400 = _T_84 ? 3'h1 : _T_399;
  wire [2:0] _T_401 = _T_82 ? 3'h0 : _T_400;
  wire [2:0] _T_402 = _T_80 ? 3'h0 : _T_401;
  wire [2:0] _T_403 = _T_78 ? 3'h0 : _T_402;
  wire [2:0] _T_404 = _T_76 ? 3'h0 : _T_403;
  wire [2:0] _T_405 = _T_74 ? 3'h0 : _T_404;
  wire [2:0] _T_406 = _T_72 ? 3'h0 : _T_405;
  wire [2:0] _T_407 = _T_70 ? 3'h0 : _T_406;
  wire [2:0] _T_408 = _T_68 ? 3'h0 : _T_407;
  wire [2:0] _T_409 = _T_66 ? 3'h0 : _T_408;
  wire [2:0] _T_410 = _T_64 ? 3'h0 : _T_409;
  wire [2:0] _T_411 = _T_62 ? 3'h0 : _T_410;
  wire [2:0] _T_412 = _T_60 ? 3'h0 : _T_411;
  wire [2:0] _T_413 = _T_58 ? 3'h0 : _T_412;
  wire [2:0] _T_414 = _T_56 ? 3'h0 : _T_413;
  wire [2:0] _T_415 = _T_54 ? 3'h0 : _T_414;
  wire [2:0] _T_416 = _T_52 ? 3'h0 : _T_415;
  wire [2:0] _T_417 = _T_50 ? 3'h0 : _T_416;
  wire [2:0] _T_418 = _T_48 ? 3'h0 : _T_417;
  wire [2:0] _T_419 = _T_46 ? 3'h0 : _T_418;
  wire [2:0] _T_420 = _T_44 ? 3'h0 : _T_419;
  wire [2:0] _T_421 = _T_42 ? 3'h0 : _T_420;
  wire [2:0] _T_422 = _T_40 ? 3'h0 : _T_421;
  wire [2:0] op2Sel = _T_38 ? 3'h0 : _T_422;
  wire [3:0] OFF26_hi_hi = inst[9] ? 4'hf : 4'h0;
  wire [9:0] OFF26_hi_lo = inst[9:0];
  wire [15:0] OFF26_lo_hi = inst[25:10];
  wire [31:0] OFF26 = {OFF26_hi_hi,OFF26_hi_lo,OFF26_lo_hi,2'h0};
  wire [19:0] UI20_hi = inst[24:5];
  wire [31:0] UI20 = {UI20_hi,12'h0};
  wire [13:0] OFF16_hi_hi = inst[25] ? 14'h3fff : 14'h0;
  wire [31:0] OFF16 = {OFF16_hi_hi,OFF26_lo_hi,2'h0};
  wire [17:0] SI14_hi = inst[23] ? 18'h3ffff : 18'h0;
  wire [13:0] SI14_lo = inst[23:10];
  wire [31:0] SI14 = {SI14_hi,SI14_lo};
  wire [19:0] SI12_hi = inst[21] ? 20'hfffff : 20'h0;
  wire [11:0] SI12_lo = inst[21:10];
  wire [31:0] SI12 = {SI12_hi,SI12_lo};
  wire [31:0] _aluOp2_WIRE_2 = {{20'd0}, SI12_lo};
  wire [4:0] k = inst[14:10];
  wire [31:0] _aluOp2_WIRE_1 = {{27'd0}, k};
  wire  _T_776 = _T_100 ? 1'h0 : _T_102;
  wire  _T_777 = _T_98 ? 1'h0 : _T_776;
  wire  _T_778 = _T_96 ? 1'h0 : _T_777;
  wire  _T_779 = _T_94 ? 1'h0 : _T_778;
  wire  _T_780 = _T_92 ? 1'h0 : _T_779;
  wire  _T_781 = _T_90 ? 1'h0 : _T_780;
  wire  _T_782 = _T_88 ? 1'h0 : _T_781;
  wire  _T_783 = _T_86 ? 1'h0 : _T_782;
  wire  _T_784 = _T_84 ? 1'h0 : _T_783;
  wire  _T_785 = _T_82 ? 1'h0 : _T_784;
  wire  _T_786 = _T_80 ? 1'h0 : _T_785;
  wire  _T_787 = _T_78 ? 1'h0 : _T_786;
  wire  _T_788 = _T_76 ? 1'h0 : _T_787;
  wire  _T_789 = _T_74 ? 1'h0 : _T_788;
  wire  _T_790 = _T_72 ? 1'h0 : _T_789;
  wire  _T_791 = _T_70 ? 1'h0 : _T_790;
  wire  _T_792 = _T_68 ? 1'h0 : _T_791;
  wire  _T_793 = _T_66 ? 1'h0 : _T_792;
  wire  _T_794 = _T_64 ? 1'h0 : _T_793;
  wire  _T_795 = _T_62 ? 1'h0 : _T_794;
  wire  _T_796 = _T_60 ? 1'h0 : _T_795;
  wire  _T_797 = _T_58 ? 1'h0 : _T_796;
  wire  _T_798 = _T_56 ? 1'h0 : _T_797;
  wire  _T_799 = _T_54 ? 1'h0 : _T_798;
  wire  _T_800 = _T_52 ? 1'h0 : _T_799;
  wire  _T_801 = _T_50 ? 1'h0 : _T_800;
  wire  _T_802 = _T_48 ? 1'h0 : _T_801;
  wire  _T_803 = _T_46 ? 1'h0 : _T_802;
  wire  _T_804 = _T_44 ? 1'h0 : _T_803;
  wire  _T_805 = _T_42 ? 1'h0 : _T_804;
  wire  _T_806 = _T_40 ? 1'h0 : _T_805;
  wire  c0_4 = _T_38 ? 1'h0 : _T_806;
  wire [2:0] _T_1127 = _T_166 ? 3'h4 : 3'h0;
  wire [2:0] _T_1128 = _T_164 ? 3'h6 : _T_1127;
  wire [2:0] _T_1129 = _T_162 ? 3'h3 : _T_1128;
  wire [2:0] _T_1130 = _T_160 ? 3'h5 : _T_1129;
  wire [2:0] _T_1131 = _T_158 ? 3'h1 : _T_1130;
  wire [2:0] _T_1132 = _T_156 ? 3'h2 : _T_1131;
  wire [2:0] _T_1133 = _T_154 ? 3'h7 : _T_1132;
  wire [2:0] _T_1134 = _T_152 ? 3'h7 : _T_1133;
  wire [2:0] _T_1135 = _T_150 ? 3'h7 : _T_1134;
  wire [2:0] _T_1136 = _T_148 ? 3'h0 : _T_1135;
  wire [2:0] _T_1137 = _T_146 ? 3'h0 : _T_1136;
  wire [2:0] _T_1138 = _T_144 ? 3'h0 : _T_1137;
  wire [2:0] _T_1139 = _T_142 ? 3'h0 : _T_1138;
  wire [2:0] _T_1140 = _T_140 ? 3'h0 : _T_1139;
  wire [2:0] _T_1141 = _T_138 ? 3'h0 : _T_1140;
  wire [2:0] _T_1142 = _T_136 ? 3'h0 : _T_1141;
  wire [2:0] _T_1143 = _T_134 ? 3'h0 : _T_1142;
  wire [2:0] _T_1144 = _T_132 ? 3'h0 : _T_1143;
  wire [2:0] _T_1145 = _T_130 ? 3'h0 : _T_1144;
  wire [2:0] _T_1146 = _T_128 ? 3'h0 : _T_1145;
  wire [2:0] _T_1147 = _T_126 ? 3'h0 : _T_1146;
  wire [2:0] _T_1148 = _T_124 ? 3'h0 : _T_1147;
  wire [2:0] _T_1149 = _T_122 ? 3'h0 : _T_1148;
  wire [2:0] _T_1150 = _T_120 ? 3'h0 : _T_1149;
  wire [2:0] _T_1151 = _T_118 ? 3'h0 : _T_1150;
  wire [2:0] _T_1152 = _T_116 ? 3'h0 : _T_1151;
  wire [2:0] _T_1153 = _T_114 ? 3'h0 : _T_1152;
  wire [2:0] _T_1154 = _T_112 ? 3'h0 : _T_1153;
  wire [2:0] _T_1155 = _T_110 ? 3'h0 : _T_1154;
  wire [2:0] _T_1156 = _T_108 ? 3'h0 : _T_1155;
  wire [2:0] _T_1157 = _T_106 ? 3'h0 : _T_1156;
  wire [2:0] _T_1158 = _T_104 ? 3'h0 : _T_1157;
  wire [2:0] _T_1159 = _T_102 ? 3'h0 : _T_1158;
  wire [2:0] _T_1160 = _T_100 ? 3'h0 : _T_1159;
  wire [2:0] _T_1161 = _T_98 ? 3'h0 : _T_1160;
  wire [2:0] _T_1162 = _T_96 ? 3'h0 : _T_1161;
  wire [2:0] _T_1163 = _T_94 ? 3'h0 : _T_1162;
  wire [2:0] _T_1164 = _T_92 ? 3'h0 : _T_1163;
  wire [2:0] _T_1165 = _T_90 ? 3'h0 : _T_1164;
  wire [2:0] _T_1166 = _T_88 ? 3'h0 : _T_1165;
  wire [2:0] _T_1167 = _T_86 ? 3'h0 : _T_1166;
  wire [2:0] _T_1168 = _T_84 ? 3'h0 : _T_1167;
  wire [2:0] _T_1169 = _T_82 ? 3'h0 : _T_1168;
  wire [2:0] _T_1170 = _T_80 ? 3'h0 : _T_1169;
  wire [2:0] _T_1171 = _T_78 ? 3'h0 : _T_1170;
  wire [2:0] _T_1172 = _T_76 ? 3'h0 : _T_1171;
  wire [2:0] _T_1173 = _T_74 ? 3'h0 : _T_1172;
  wire [2:0] _T_1174 = _T_72 ? 3'h0 : _T_1173;
  wire [2:0] _T_1175 = _T_70 ? 3'h0 : _T_1174;
  wire [2:0] _T_1176 = _T_68 ? 3'h0 : _T_1175;
  wire [2:0] _T_1177 = _T_66 ? 3'h0 : _T_1176;
  wire [2:0] _T_1178 = _T_64 ? 3'h0 : _T_1177;
  wire [2:0] _T_1179 = _T_62 ? 3'h0 : _T_1178;
  wire [2:0] _T_1180 = _T_60 ? 3'h0 : _T_1179;
  wire [2:0] _T_1181 = _T_58 ? 3'h0 : _T_1180;
  wire [2:0] _T_1182 = _T_56 ? 3'h0 : _T_1181;
  wire [2:0] _T_1183 = _T_54 ? 3'h0 : _T_1182;
  wire [2:0] _T_1184 = _T_52 ? 3'h0 : _T_1183;
  wire [2:0] _T_1185 = _T_50 ? 3'h0 : _T_1184;
  wire [2:0] _T_1186 = _T_48 ? 3'h0 : _T_1185;
  wire [2:0] _T_1187 = _T_46 ? 3'h0 : _T_1186;
  wire [2:0] _T_1188 = _T_44 ? 3'h0 : _T_1187;
  wire [2:0] _T_1189 = _T_42 ? 3'h0 : _T_1188;
  wire [2:0] _T_1190 = _T_40 ? 3'h0 : _T_1189;
  wire [2:0] brType = _T_38 ? 3'h0 : _T_1190;
  wire  _kd_T_5 = ~(&c0_3[2:1]) | c0_4 | |brType;
  wire [4:0] kd = ~(&c0_3[2:1]) | c0_4 | |brType ? d : k;
  wire [31:0] rkd = kd == 5'h0 ? 32'h0 : GR_rkd_MPORT_data;
  wire [31:0] _GEN_61 = 3'h1 == op2Sel ? _aluOp2_WIRE_1 : rkd;
  wire [31:0] _GEN_62 = 3'h2 == op2Sel ? _aluOp2_WIRE_2 : _GEN_61;
  wire [31:0] _GEN_63 = 3'h3 == op2Sel ? SI12 : _GEN_62;
  wire [31:0] _GEN_64 = 3'h4 == op2Sel ? SI14 : _GEN_63;
  wire [31:0] _GEN_65 = 3'h5 == op2Sel ? OFF16 : _GEN_64;
  wire [31:0] _GEN_66 = 3'h6 == op2Sel ? UI20 : _GEN_65;
  wire [31:0] _GEN_67 = 3'h7 == op2Sel ? OFF26 : _GEN_66;
  wire [31:0] _aluOut_T_2 = aluOp1 + _GEN_67;
  wire [31:0] _aluOut_T_65 = _aluOut_T ? _aluOut_T_2 : 32'h0;
  wire  _aluOut_T_4 = func == 5'h1;
  wire [31:0] _aluOut_T_6 = aluOp1 - _GEN_67;
  wire [31:0] _aluOut_T_66 = _aluOut_T_4 ? _aluOut_T_6 : 32'h0;
  wire [31:0] _aluOut_T_84 = _aluOut_T_65 | _aluOut_T_66;
  wire  _aluOut_T_8 = func == 5'h2;
  wire [62:0] _GEN_4317 = {{31'd0}, aluOp1};
  wire [62:0] _aluOut_T_10 = _GEN_4317 << _GEN_67[4:0];
  wire [31:0] _aluOut_T_67 = _aluOut_T_8 ? _aluOut_T_10[31:0] : 32'h0;
  wire [31:0] _aluOut_T_85 = _aluOut_T_84 | _aluOut_T_67;
  wire  _aluOut_T_12 = func == 5'h3;
  wire [31:0] _aluOut_T_14 = aluOp1 >> _GEN_67[4:0];
  wire [31:0] _aluOut_T_68 = _aluOut_T_12 ? _aluOut_T_14 : 32'h0;
  wire [31:0] _aluOut_T_86 = _aluOut_T_85 | _aluOut_T_68;
  wire  _aluOut_T_16 = func == 5'h4;
  wire [31:0] aluOut_sa = ~op1Sel ? rj : PC;
  wire [31:0] _aluOut_T_19 = $signed(aluOut_sa) >>> _GEN_67[4:0];
  wire [31:0] _aluOut_T_69 = _aluOut_T_16 ? _aluOut_T_19 : 32'h0;
  wire [31:0] _aluOut_T_87 = _aluOut_T_86 | _aluOut_T_69;
  wire  _aluOut_T_21 = func == 5'h5;
  wire [31:0] _aluOut_T_22 = aluOp1 & _GEN_67;
  wire [31:0] _aluOut_T_70 = _aluOut_T_21 ? _aluOut_T_22 : 32'h0;
  wire [31:0] _aluOut_T_88 = _aluOut_T_87 | _aluOut_T_70;
  wire  _aluOut_T_24 = func == 5'h6;
  wire [31:0] _aluOut_T_25 = aluOp1 | _GEN_67;
  wire [31:0] _aluOut_T_71 = _aluOut_T_24 ? _aluOut_T_25 : 32'h0;
  wire [31:0] _aluOut_T_89 = _aluOut_T_88 | _aluOut_T_71;
  wire  _aluOut_T_27 = func == 5'h7;
  wire [31:0] _aluOut_T_29 = ~_aluOut_T_25;
  wire [31:0] _aluOut_T_72 = _aluOut_T_27 ? _aluOut_T_29 : 32'h0;
  wire [31:0] _aluOut_T_90 = _aluOut_T_89 | _aluOut_T_72;
  wire  _aluOut_T_31 = func == 5'h8;
  wire [31:0] _aluOut_T_32 = aluOp1 ^ _GEN_67;
  wire [31:0] _aluOut_T_73 = _aluOut_T_31 ? _aluOut_T_32 : 32'h0;
  wire [31:0] _aluOut_T_91 = _aluOut_T_90 | _aluOut_T_73;
  wire  _aluOut_T_34 = func == 5'h9;
  wire [31:0] aluOut_sb = 3'h7 == op2Sel ? OFF26 : _GEN_66;
  wire  _aluOut_T_35 = $signed(aluOut_sa) < $signed(aluOut_sb);
  wire  _aluOut_T_74 = _aluOut_T_34 & _aluOut_T_35;
  wire [31:0] _GEN_4318 = {{31'd0}, _aluOut_T_74};
  wire [31:0] _aluOut_T_92 = _aluOut_T_91 | _GEN_4318;
  wire  _aluOut_T_36 = func == 5'ha;
  wire  _aluOut_T_37 = aluOp1 < _GEN_67;
  wire  _aluOut_T_75 = _aluOut_T_36 & _aluOut_T_37;
  wire [31:0] _GEN_4319 = {{31'd0}, _aluOut_T_75};
  wire [31:0] _aluOut_T_93 = _aluOut_T_92 | _GEN_4319;
  wire  _aluOut_T_38 = func == 5'hb;
  wire [31:0] _aluOut_T_76 = _aluOut_T_38 ? _GEN_67 : 32'h0;
  wire [31:0] _aluOut_T_94 = _aluOut_T_93 | _aluOut_T_76;
  wire  _aluOut_T_40 = func == 5'hc;
  wire [63:0] _aluOut_T_42 = $signed(aluOut_sa) * $signed(aluOut_sb);
  wire [31:0] _aluOut_T_77 = _aluOut_T_40 ? _aluOut_T_42[31:0] : 32'h0;
  wire [31:0] _aluOut_T_95 = _aluOut_T_94 | _aluOut_T_77;
  wire  _aluOut_T_44 = func == 5'hd;
  wire [31:0] _aluOut_T_78 = _aluOut_T_44 ? _aluOut_T_42[63:32] : 32'h0;
  wire [31:0] _aluOut_T_96 = _aluOut_T_95 | _aluOut_T_78;
  wire  _aluOut_T_48 = func == 5'he;
  wire [63:0] _aluOut_T_49 = aluOp1 * _GEN_67;
  wire [31:0] _aluOut_T_79 = _aluOut_T_48 ? _aluOut_T_49[63:32] : 32'h0;
  wire [31:0] _aluOut_T_97 = _aluOut_T_96 | _aluOut_T_79;
  wire  _aluOut_T_51 = func == 5'hf;
  wire [31:0] _aluOut_T_53 = $signed(aluOut_sa) % $signed(aluOut_sb);
  wire [31:0] _aluOut_T_80 = _aluOut_T_51 ? _aluOut_T_53 : 32'h0;
  wire [31:0] _aluOut_T_98 = _aluOut_T_97 | _aluOut_T_80;
  wire  _aluOut_T_55 = func == 5'h10;
  wire [32:0] _aluOut_T_57 = $signed(aluOut_sa) / $signed(aluOut_sb);
  wire [31:0] _aluOut_T_81 = _aluOut_T_55 ? _aluOut_T_57[31:0] : 32'h0;
  wire [31:0] _aluOut_T_99 = _aluOut_T_98 | _aluOut_T_81;
  wire  _aluOut_T_59 = func == 5'h11;
  wire [31:0] _GEN_9 = aluOp1 % _GEN_67;
  wire [31:0] _aluOut_T_60 = _GEN_9[31:0];
  wire [31:0] _aluOut_T_82 = _aluOut_T_59 ? _aluOut_T_60 : 32'h0;
  wire [31:0] _aluOut_T_100 = _aluOut_T_99 | _aluOut_T_82;
  wire  _aluOut_T_62 = func == 5'h12;
  wire [31:0] _aluOut_T_63 = aluOp1 / _GEN_67;
  wire [31:0] _aluOut_T_83 = _aluOut_T_62 ? _aluOut_T_63 : 32'h0;
  wire [31:0] aluOut = _aluOut_T_100 | _aluOut_T_83;
  wire  memALE = aluOut[0] & c0_3[2:1] == 2'h1 | |aluOut[1:0] & c0_3[2:1] == 2'h2;
  wire  memADEM = aluOut[31] & _T_32;
  wire  _EXVA_T = c0_3 != 3'h7;
  wire [31:0] _EXVA_T_4 = _EXVA_T ? aluOut : 32'h0;
  wire [2:0] _T_961 = _T_114 ? 3'h5 : 3'h0;
  wire [2:0] _T_962 = _T_112 ? 3'h4 : _T_961;
  wire [2:0] _T_963 = _T_110 ? 3'h3 : _T_962;
  wire [2:0] _T_964 = _T_108 ? 3'h2 : _T_963;
  wire [2:0] _T_965 = _T_106 ? 3'h1 : _T_964;
  wire [2:0] _T_966 = _T_104 ? 3'h0 : _T_965;
  wire [2:0] _T_967 = _T_102 ? 3'h0 : _T_966;
  wire [2:0] _T_968 = _T_100 ? 3'h0 : _T_967;
  wire [2:0] _T_969 = _T_98 ? 3'h0 : _T_968;
  wire [2:0] _T_970 = _T_96 ? 3'h0 : _T_969;
  wire [2:0] _T_971 = _T_94 ? 3'h0 : _T_970;
  wire [2:0] _T_972 = _T_92 ? 3'h0 : _T_971;
  wire [2:0] _T_973 = _T_90 ? 3'h0 : _T_972;
  wire [2:0] _T_974 = _T_88 ? 3'h0 : _T_973;
  wire [2:0] _T_975 = _T_86 ? 3'h0 : _T_974;
  wire [2:0] _T_976 = _T_84 ? 3'h0 : _T_975;
  wire [2:0] _T_977 = _T_82 ? 3'h0 : _T_976;
  wire [2:0] _T_978 = _T_80 ? 3'h0 : _T_977;
  wire [2:0] _T_979 = _T_78 ? 3'h0 : _T_978;
  wire [2:0] _T_980 = _T_76 ? 3'h0 : _T_979;
  wire [2:0] _T_981 = _T_74 ? 3'h0 : _T_980;
  wire [2:0] _T_982 = _T_72 ? 3'h0 : _T_981;
  wire [2:0] _T_983 = _T_70 ? 3'h0 : _T_982;
  wire [2:0] _T_984 = _T_68 ? 3'h0 : _T_983;
  wire [2:0] _T_985 = _T_66 ? 3'h0 : _T_984;
  wire [2:0] _T_986 = _T_64 ? 3'h0 : _T_985;
  wire [2:0] _T_987 = _T_62 ? 3'h0 : _T_986;
  wire [2:0] _T_988 = _T_60 ? 3'h0 : _T_987;
  wire [2:0] _T_989 = _T_58 ? 3'h0 : _T_988;
  wire [2:0] _T_990 = _T_56 ? 3'h0 : _T_989;
  wire [2:0] _T_991 = _T_54 ? 3'h0 : _T_990;
  wire [2:0] _T_992 = _T_52 ? 3'h0 : _T_991;
  wire [2:0] _T_993 = _T_50 ? 3'h0 : _T_992;
  wire [2:0] _T_994 = _T_48 ? 3'h0 : _T_993;
  wire [2:0] _T_995 = _T_46 ? 3'h0 : _T_994;
  wire [2:0] _T_996 = _T_44 ? 3'h0 : _T_995;
  wire [2:0] _T_997 = _T_42 ? 3'h0 : _T_996;
  wire [2:0] _T_998 = _T_40 ? 3'h0 : _T_997;
  wire [2:0] c0_7 = _T_38 ? 3'h0 : _T_998;
  wire  _EXVA_T_1 = c0_7 == 3'h1;
  wire [31:0] _EXVA_T_2 = {csrs_9_VPPN,13'h0};
  wire [31:0] _EXVA_T_5 = _EXVA_T_1 ? _EXVA_T_2 : 32'h0;
  wire [31:0] _EXVA_T_7 = _EXVA_T_4 | _EXVA_T_5;
  wire  _EXVA_T_3 = c0_7 == 3'h5;
  wire [31:0] _EXVA_T_6 = _EXVA_T_3 ? rkd : 32'h0;
  wire [31:0] EXVA = _EXVA_T_7 | _EXVA_T_6;
  wire  vaMatch_0_1 = tlb_0_VPPN[18:10] == EXVA[31:23] & (tlb_0_PS == 6'h16 | tlb_0_VPPN[9:0] == EXVA[22:13]);
  wire [9:0] EXASID = _EXVA_T_3 ? rj[9:0] : asid_ASID;
  wire  asidMatch_0_1 = tlb_0_ASID == EXASID;
  wire  tlbHit_0_1 = tlb_0_E & vaMatch_0_1 & (tlb_0_G | asidMatch_0_1);
  wire  vaMatch_1_1 = tlb_1_VPPN[18:10] == EXVA[31:23] & (tlb_1_PS == 6'h16 | tlb_1_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_1_1 = tlb_1_ASID == EXASID;
  wire  tlbHit_1_1 = tlb_1_E & vaMatch_1_1 & (tlb_1_G | asidMatch_1_1);
  wire  vaMatch_2_1 = tlb_2_VPPN[18:10] == EXVA[31:23] & (tlb_2_PS == 6'h16 | tlb_2_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_2_1 = tlb_2_ASID == EXASID;
  wire  tlbHit_2_1 = tlb_2_E & vaMatch_2_1 & (tlb_2_G | asidMatch_2_1);
  wire  vaMatch_3_1 = tlb_3_VPPN[18:10] == EXVA[31:23] & (tlb_3_PS == 6'h16 | tlb_3_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_3_1 = tlb_3_ASID == EXASID;
  wire  tlbHit_3_1 = tlb_3_E & vaMatch_3_1 & (tlb_3_G | asidMatch_3_1);
  wire  vaMatch_4_1 = tlb_4_VPPN[18:10] == EXVA[31:23] & (tlb_4_PS == 6'h16 | tlb_4_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_4_1 = tlb_4_ASID == EXASID;
  wire  tlbHit_4_1 = tlb_4_E & vaMatch_4_1 & (tlb_4_G | asidMatch_4_1);
  wire  vaMatch_5_1 = tlb_5_VPPN[18:10] == EXVA[31:23] & (tlb_5_PS == 6'h16 | tlb_5_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_5_1 = tlb_5_ASID == EXASID;
  wire  tlbHit_5_1 = tlb_5_E & vaMatch_5_1 & (tlb_5_G | asidMatch_5_1);
  wire  vaMatch_6_1 = tlb_6_VPPN[18:10] == EXVA[31:23] & (tlb_6_PS == 6'h16 | tlb_6_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_6_1 = tlb_6_ASID == EXASID;
  wire  tlbHit_6_1 = tlb_6_E & vaMatch_6_1 & (tlb_6_G | asidMatch_6_1);
  wire  vaMatch_7_1 = tlb_7_VPPN[18:10] == EXVA[31:23] & (tlb_7_PS == 6'h16 | tlb_7_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_7_1 = tlb_7_ASID == EXASID;
  wire  tlbHit_7_1 = tlb_7_E & vaMatch_7_1 & (tlb_7_G | asidMatch_7_1);
  wire  vaMatch_8_1 = tlb_8_VPPN[18:10] == EXVA[31:23] & (tlb_8_PS == 6'h16 | tlb_8_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_8_1 = tlb_8_ASID == EXASID;
  wire  tlbHit_8_1 = tlb_8_E & vaMatch_8_1 & (tlb_8_G | asidMatch_8_1);
  wire  vaMatch_9_1 = tlb_9_VPPN[18:10] == EXVA[31:23] & (tlb_9_PS == 6'h16 | tlb_9_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_9_1 = tlb_9_ASID == EXASID;
  wire  tlbHit_9_1 = tlb_9_E & vaMatch_9_1 & (tlb_9_G | asidMatch_9_1);
  wire  vaMatch_10_1 = tlb_10_VPPN[18:10] == EXVA[31:23] & (tlb_10_PS == 6'h16 | tlb_10_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_10_1 = tlb_10_ASID == EXASID;
  wire  tlbHit_10_1 = tlb_10_E & vaMatch_10_1 & (tlb_10_G | asidMatch_10_1);
  wire  vaMatch_11_1 = tlb_11_VPPN[18:10] == EXVA[31:23] & (tlb_11_PS == 6'h16 | tlb_11_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_11_1 = tlb_11_ASID == EXASID;
  wire  tlbHit_11_1 = tlb_11_E & vaMatch_11_1 & (tlb_11_G | asidMatch_11_1);
  wire  vaMatch_12_1 = tlb_12_VPPN[18:10] == EXVA[31:23] & (tlb_12_PS == 6'h16 | tlb_12_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_12_1 = tlb_12_ASID == EXASID;
  wire  tlbHit_12_1 = tlb_12_E & vaMatch_12_1 & (tlb_12_G | asidMatch_12_1);
  wire  vaMatch_13_1 = tlb_13_VPPN[18:10] == EXVA[31:23] & (tlb_13_PS == 6'h16 | tlb_13_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_13_1 = tlb_13_ASID == EXASID;
  wire  tlbHit_13_1 = tlb_13_E & vaMatch_13_1 & (tlb_13_G | asidMatch_13_1);
  wire  vaMatch_14_1 = tlb_14_VPPN[18:10] == EXVA[31:23] & (tlb_14_PS == 6'h16 | tlb_14_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_14_1 = tlb_14_ASID == EXASID;
  wire  tlbHit_14_1 = tlb_14_E & vaMatch_14_1 & (tlb_14_G | asidMatch_14_1);
  wire  vaMatch_15_1 = tlb_15_VPPN[18:10] == EXVA[31:23] & (tlb_15_PS == 6'h16 | tlb_15_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_15_1 = tlb_15_ASID == EXASID;
  wire  tlbHit_15_1 = tlb_15_E & vaMatch_15_1 & (tlb_15_G | asidMatch_15_1);
  wire  vaMatch_16_1 = tlb_16_VPPN[18:10] == EXVA[31:23] & (tlb_16_PS == 6'h16 | tlb_16_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_16_1 = tlb_16_ASID == EXASID;
  wire  tlbHit_16_1 = tlb_16_E & vaMatch_16_1 & (tlb_16_G | asidMatch_16_1);
  wire  vaMatch_17_1 = tlb_17_VPPN[18:10] == EXVA[31:23] & (tlb_17_PS == 6'h16 | tlb_17_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_17_1 = tlb_17_ASID == EXASID;
  wire  tlbHit_17_1 = tlb_17_E & vaMatch_17_1 & (tlb_17_G | asidMatch_17_1);
  wire  vaMatch_18_1 = tlb_18_VPPN[18:10] == EXVA[31:23] & (tlb_18_PS == 6'h16 | tlb_18_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_18_1 = tlb_18_ASID == EXASID;
  wire  tlbHit_18_1 = tlb_18_E & vaMatch_18_1 & (tlb_18_G | asidMatch_18_1);
  wire  vaMatch_19_1 = tlb_19_VPPN[18:10] == EXVA[31:23] & (tlb_19_PS == 6'h16 | tlb_19_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_19_1 = tlb_19_ASID == EXASID;
  wire  tlbHit_19_1 = tlb_19_E & vaMatch_19_1 & (tlb_19_G | asidMatch_19_1);
  wire  vaMatch_20_1 = tlb_20_VPPN[18:10] == EXVA[31:23] & (tlb_20_PS == 6'h16 | tlb_20_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_20_1 = tlb_20_ASID == EXASID;
  wire  tlbHit_20_1 = tlb_20_E & vaMatch_20_1 & (tlb_20_G | asidMatch_20_1);
  wire  vaMatch_21_1 = tlb_21_VPPN[18:10] == EXVA[31:23] & (tlb_21_PS == 6'h16 | tlb_21_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_21_1 = tlb_21_ASID == EXASID;
  wire  tlbHit_21_1 = tlb_21_E & vaMatch_21_1 & (tlb_21_G | asidMatch_21_1);
  wire  vaMatch_22_1 = tlb_22_VPPN[18:10] == EXVA[31:23] & (tlb_22_PS == 6'h16 | tlb_22_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_22_1 = tlb_22_ASID == EXASID;
  wire  tlbHit_22_1 = tlb_22_E & vaMatch_22_1 & (tlb_22_G | asidMatch_22_1);
  wire  vaMatch_23_1 = tlb_23_VPPN[18:10] == EXVA[31:23] & (tlb_23_PS == 6'h16 | tlb_23_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_23_1 = tlb_23_ASID == EXASID;
  wire  tlbHit_23_1 = tlb_23_E & vaMatch_23_1 & (tlb_23_G | asidMatch_23_1);
  wire  vaMatch_24_1 = tlb_24_VPPN[18:10] == EXVA[31:23] & (tlb_24_PS == 6'h16 | tlb_24_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_24_1 = tlb_24_ASID == EXASID;
  wire  tlbHit_24_1 = tlb_24_E & vaMatch_24_1 & (tlb_24_G | asidMatch_24_1);
  wire  vaMatch_25_1 = tlb_25_VPPN[18:10] == EXVA[31:23] & (tlb_25_PS == 6'h16 | tlb_25_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_25_1 = tlb_25_ASID == EXASID;
  wire  tlbHit_25_1 = tlb_25_E & vaMatch_25_1 & (tlb_25_G | asidMatch_25_1);
  wire  vaMatch_26_1 = tlb_26_VPPN[18:10] == EXVA[31:23] & (tlb_26_PS == 6'h16 | tlb_26_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_26_1 = tlb_26_ASID == EXASID;
  wire  tlbHit_26_1 = tlb_26_E & vaMatch_26_1 & (tlb_26_G | asidMatch_26_1);
  wire  vaMatch_27_1 = tlb_27_VPPN[18:10] == EXVA[31:23] & (tlb_27_PS == 6'h16 | tlb_27_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_27_1 = tlb_27_ASID == EXASID;
  wire  tlbHit_27_1 = tlb_27_E & vaMatch_27_1 & (tlb_27_G | asidMatch_27_1);
  wire  vaMatch_28_1 = tlb_28_VPPN[18:10] == EXVA[31:23] & (tlb_28_PS == 6'h16 | tlb_28_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_28_1 = tlb_28_ASID == EXASID;
  wire  tlbHit_28_1 = tlb_28_E & vaMatch_28_1 & (tlb_28_G | asidMatch_28_1);
  wire  vaMatch_29_1 = tlb_29_VPPN[18:10] == EXVA[31:23] & (tlb_29_PS == 6'h16 | tlb_29_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_29_1 = tlb_29_ASID == EXASID;
  wire  tlbHit_29_1 = tlb_29_E & vaMatch_29_1 & (tlb_29_G | asidMatch_29_1);
  wire  vaMatch_30_1 = tlb_30_VPPN[18:10] == EXVA[31:23] & (tlb_30_PS == 6'h16 | tlb_30_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_30_1 = tlb_30_ASID == EXASID;
  wire  tlbHit_30_1 = tlb_30_E & vaMatch_30_1 & (tlb_30_G | asidMatch_30_1);
  wire  _miss_T_61 = tlbHit_0_1 | tlbHit_1_1 | tlbHit_2_1 | tlbHit_3_1 | tlbHit_4_1 | tlbHit_5_1 | tlbHit_6_1 |
    tlbHit_7_1 | tlbHit_8_1 | tlbHit_9_1 | tlbHit_10_1 | tlbHit_11_1 | tlbHit_12_1 | tlbHit_13_1 | tlbHit_14_1 |
    tlbHit_15_1 | tlbHit_16_1 | tlbHit_17_1 | tlbHit_18_1 | tlbHit_19_1 | tlbHit_20_1 | tlbHit_21_1 | tlbHit_22_1 |
    tlbHit_23_1 | tlbHit_24_1 | tlbHit_25_1 | tlbHit_26_1 | tlbHit_27_1 | tlbHit_28_1 | tlbHit_29_1 | tlbHit_30_1;
  wire  vaMatch_31_1 = tlb_31_VPPN[18:10] == EXVA[31:23] & (tlb_31_PS == 6'h16 | tlb_31_VPPN[9:0] == EXVA[22:13]);
  wire  asidMatch_31_1 = tlb_31_ASID == EXASID;
  wire  tlbHit_31_1 = tlb_31_E & vaMatch_31_1 & (tlb_31_G | asidMatch_31_1);
  wire  _miss_T_62 = _miss_T_61 | tlbHit_31_1;
  wire  _GEN_70 = EXVA[31:29] == csrs_28_VSEG & (csrs_28_PLV0 & _T_11 | csrs_28_PLV3 & _T_13) ? 1'h0 : ~(_miss_T_61 |
    tlbHit_31_1);
  wire  miss_1 = EXVA[31:29] == csrs_27_VSEG & (csrs_27_PLV0 & crmd_PLV == 2'h0 | csrs_27_PLV3 & crmd_PLV == 2'h3) ? 1'h0
     : _GEN_70;
  wire  _T_1267 = _T_142 ? 1'h0 : _T_144;
  wire  _T_1268 = _T_140 ? 1'h0 : _T_1267;
  wire  _T_1269 = _T_138 ? 1'h0 : _T_1268;
  wire  _T_1270 = _T_136 ? 1'h0 : _T_1269;
  wire  _T_1271 = _T_134 ? 1'h0 : _T_1270;
  wire  _T_1272 = _T_132 ? 1'h0 : _T_1271;
  wire  _T_1273 = _T_130 ? 1'h0 : _T_1272;
  wire  _T_1274 = _T_128 ? 1'h0 : _T_1273;
  wire  _T_1275 = _T_126 ? 1'h0 : _T_1274;
  wire  _T_1276 = _T_124 ? 1'h0 : _T_1275;
  wire  _T_1277 = _T_122 ? 1'h0 : _T_1276;
  wire  _T_1278 = _T_120 ? 1'h0 : _T_1277;
  wire  _T_1279 = _T_118 ? 1'h0 : _T_1278;
  wire  _T_1280 = _T_116 ? 1'h0 : _T_1279;
  wire  _T_1281 = _T_114 ? 1'h0 : _T_1280;
  wire  _T_1282 = _T_112 ? 1'h0 : _T_1281;
  wire  _T_1283 = _T_110 ? 1'h0 : _T_1282;
  wire  _T_1284 = _T_108 ? 1'h0 : _T_1283;
  wire  _T_1285 = _T_106 ? 1'h0 : _T_1284;
  wire  _T_1286 = _T_104 ? 1'h0 : _T_1285;
  wire  _T_1287 = _T_102 ? 1'h0 : _T_1286;
  wire  _T_1288 = _T_100 ? 1'h0 : _T_1287;
  wire  _T_1289 = _T_98 ? 1'h0 : _T_1288;
  wire  _T_1290 = _T_96 ? 1'h0 : _T_1289;
  wire  _T_1291 = _T_94 ? 1'h0 : _T_1290;
  wire  _T_1292 = _T_92 ? 1'h0 : _T_1291;
  wire  _T_1293 = _T_90 ? 1'h0 : _T_1292;
  wire  _T_1294 = _T_88 ? 1'h0 : _T_1293;
  wire  _T_1295 = _T_86 ? 1'h0 : _T_1294;
  wire  _T_1296 = _T_84 ? 1'h0 : _T_1295;
  wire  _T_1297 = _T_82 ? 1'h0 : _T_1296;
  wire  _T_1298 = _T_80 ? 1'h0 : _T_1297;
  wire  _T_1299 = _T_78 ? 1'h0 : _T_1298;
  wire  _T_1300 = _T_76 ? 1'h0 : _T_1299;
  wire  _T_1301 = _T_74 ? 1'h0 : _T_1300;
  wire  _T_1302 = _T_72 ? 1'h0 : _T_1301;
  wire  _T_1303 = _T_70 ? 1'h0 : _T_1302;
  wire  _T_1304 = _T_68 ? 1'h0 : _T_1303;
  wire  _T_1305 = _T_66 ? 1'h0 : _T_1304;
  wire  _T_1306 = _T_64 ? 1'h0 : _T_1305;
  wire  _T_1307 = _T_62 ? 1'h0 : _T_1306;
  wire  _T_1308 = _T_60 ? 1'h0 : _T_1307;
  wire  _T_1309 = _T_58 ? 1'h0 : _T_1308;
  wire  _T_1310 = _T_56 ? 1'h0 : _T_1309;
  wire  _T_1311 = _T_54 ? 1'h0 : _T_1310;
  wire  _T_1312 = _T_52 ? 1'h0 : _T_1311;
  wire  _T_1313 = _T_50 ? 1'h0 : _T_1312;
  wire  _T_1314 = _T_48 ? 1'h0 : _T_1313;
  wire  _T_1315 = _T_46 ? 1'h0 : _T_1314;
  wire  _T_1316 = _T_44 ? 1'h0 : _T_1315;
  wire  _T_1317 = _T_42 ? 1'h0 : _T_1316;
  wire  _T_1318 = _T_40 ? 1'h0 : _T_1317;
  wire  c0_12 = _T_38 ? 1'h0 : _T_1318;
  wire  _lo_T_2 = ~c0_12;
  wire  _GEN_100 = miss_1 ? ~c0_12 : _GEN_45;
  wire  _GEN_108 = crmd_DA ? _GEN_45 : _GEN_100;
  wire  _GEN_116 = memADEM ? _GEN_45 : _GEN_108;
  wire  _GEN_125 = memALE ? _GEN_45 : _GEN_116;
  wire  _GEN_134 = c0_3 == 3'h7 | c0_11 & d[4:3] != 2'h2 ? _GEN_45 : _GEN_125;
  wire  _GEN_148 = ID_OK ? _GEN_134 : _GEN_45;
  wire  TLBR = dStallReg ? _GEN_45 : _GEN_148;
  wire  _GEN_53 = IF_OK & ~iStall & break_;
  wire  BRK = dStallReg ? 1'h0 : _GEN_53;
  wire  _T_1443 = 3'h1 == c0_7;
  wire  _GEN_54 = IF_OK & ~iStall & ~instV;
  wire  _GEN_59 = dStallReg ? 1'h0 : _GEN_54;
  wire  _T_1475 = 3'h2 == c0_7;
  wire  _T_1476 = 3'h3 == c0_7;
  wire  _T_1477 = 3'h4 == c0_7;
  wire  _T_1479 = 3'h5 == c0_7;
  wire  inv_op_0 = d == 5'h0 | d == 5'h1;
  wire  inv_op_1 = d == 5'h2;
  wire  inv_op_2 = d == 5'h3;
  wire  inv_op_3 = d == 5'h4;
  wire  inv_op_4 = d == 5'h5;
  wire  inv_op_5 = d == 5'h6;
  wire  _GEN_1777 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? _GEN_59 : 1'h1;
  wire  _GEN_1810 = _T_1479 ? _GEN_1777 : _GEN_59;
  wire  _GEN_2291 = _T_1477 ? _GEN_59 : _GEN_1810;
  wire  _GEN_2772 = _T_1476 ? _GEN_59 : _GEN_2291;
  wire  _GEN_3269 = _T_1475 ? _GEN_59 : _GEN_2772;
  wire  _GEN_3767 = _T_1443 ? _GEN_59 : _GEN_3269;
  wire  INE = ID_OK ? _GEN_3767 : _GEN_59;
  wire  _GEN_122 = memALE & _lo_T_2;
  wire  _GEN_132 = c0_3 == 3'h7 | c0_11 & d[4:3] != 2'h2 ? 1'h0 : _GEN_122;
  wire  _GEN_146 = ID_OK & _GEN_132;
  wire  ALE = dStallReg ? 1'h0 : _GEN_146;
  wire  _GEN_52 = IF_OK & ~iStall & c0_6;
  wire  SYS = dStallReg ? 1'h0 : _GEN_52;
  wire [7:0] excp_lo = {ALE,SYS,BRK,INE,2'h0,1'h0,TLBR};
  wire  _GEN_38 = ~INT & ~idle & _T_34;
  wire  ADEF = dStallReg | iStallReg ? 1'h0 : _GEN_38;
  wire  _GEN_114 = memADEM & _lo_T_2;
  wire  _GEN_123 = memALE ? 1'h0 : _GEN_114;
  wire  _GEN_133 = c0_3 == 3'h7 | c0_11 & d[4:3] != 2'h2 ? 1'h0 : _GEN_123;
  wire  _GEN_147 = ID_OK & _GEN_133;
  wire  ADEM = dStallReg ? 1'h0 : _GEN_147;
  wire [5:0] _foundTLB_T_1764 = tlbHit_0_1 ? tlb_0_PS : 6'h0;
  wire [5:0] _foundTLB_T_1765 = tlbHit_1_1 ? tlb_1_PS : 6'h0;
  wire [5:0] _foundTLB_T_1796 = _foundTLB_T_1764 | _foundTLB_T_1765;
  wire [5:0] _foundTLB_T_1766 = tlbHit_2_1 ? tlb_2_PS : 6'h0;
  wire [5:0] _foundTLB_T_1797 = _foundTLB_T_1796 | _foundTLB_T_1766;
  wire [5:0] _foundTLB_T_1767 = tlbHit_3_1 ? tlb_3_PS : 6'h0;
  wire [5:0] _foundTLB_T_1798 = _foundTLB_T_1797 | _foundTLB_T_1767;
  wire [5:0] _foundTLB_T_1768 = tlbHit_4_1 ? tlb_4_PS : 6'h0;
  wire [5:0] _foundTLB_T_1799 = _foundTLB_T_1798 | _foundTLB_T_1768;
  wire [5:0] _foundTLB_T_1769 = tlbHit_5_1 ? tlb_5_PS : 6'h0;
  wire [5:0] _foundTLB_T_1800 = _foundTLB_T_1799 | _foundTLB_T_1769;
  wire [5:0] _foundTLB_T_1770 = tlbHit_6_1 ? tlb_6_PS : 6'h0;
  wire [5:0] _foundTLB_T_1801 = _foundTLB_T_1800 | _foundTLB_T_1770;
  wire [5:0] _foundTLB_T_1771 = tlbHit_7_1 ? tlb_7_PS : 6'h0;
  wire [5:0] _foundTLB_T_1802 = _foundTLB_T_1801 | _foundTLB_T_1771;
  wire [5:0] _foundTLB_T_1772 = tlbHit_8_1 ? tlb_8_PS : 6'h0;
  wire [5:0] _foundTLB_T_1803 = _foundTLB_T_1802 | _foundTLB_T_1772;
  wire [5:0] _foundTLB_T_1773 = tlbHit_9_1 ? tlb_9_PS : 6'h0;
  wire [5:0] _foundTLB_T_1804 = _foundTLB_T_1803 | _foundTLB_T_1773;
  wire [5:0] _foundTLB_T_1774 = tlbHit_10_1 ? tlb_10_PS : 6'h0;
  wire [5:0] _foundTLB_T_1805 = _foundTLB_T_1804 | _foundTLB_T_1774;
  wire [5:0] _foundTLB_T_1775 = tlbHit_11_1 ? tlb_11_PS : 6'h0;
  wire [5:0] _foundTLB_T_1806 = _foundTLB_T_1805 | _foundTLB_T_1775;
  wire [5:0] _foundTLB_T_1776 = tlbHit_12_1 ? tlb_12_PS : 6'h0;
  wire [5:0] _foundTLB_T_1807 = _foundTLB_T_1806 | _foundTLB_T_1776;
  wire [5:0] _foundTLB_T_1777 = tlbHit_13_1 ? tlb_13_PS : 6'h0;
  wire [5:0] _foundTLB_T_1808 = _foundTLB_T_1807 | _foundTLB_T_1777;
  wire [5:0] _foundTLB_T_1778 = tlbHit_14_1 ? tlb_14_PS : 6'h0;
  wire [5:0] _foundTLB_T_1809 = _foundTLB_T_1808 | _foundTLB_T_1778;
  wire [5:0] _foundTLB_T_1779 = tlbHit_15_1 ? tlb_15_PS : 6'h0;
  wire [5:0] _foundTLB_T_1810 = _foundTLB_T_1809 | _foundTLB_T_1779;
  wire [5:0] _foundTLB_T_1780 = tlbHit_16_1 ? tlb_16_PS : 6'h0;
  wire [5:0] _foundTLB_T_1811 = _foundTLB_T_1810 | _foundTLB_T_1780;
  wire [5:0] _foundTLB_T_1781 = tlbHit_17_1 ? tlb_17_PS : 6'h0;
  wire [5:0] _foundTLB_T_1812 = _foundTLB_T_1811 | _foundTLB_T_1781;
  wire [5:0] _foundTLB_T_1782 = tlbHit_18_1 ? tlb_18_PS : 6'h0;
  wire [5:0] _foundTLB_T_1813 = _foundTLB_T_1812 | _foundTLB_T_1782;
  wire [5:0] _foundTLB_T_1783 = tlbHit_19_1 ? tlb_19_PS : 6'h0;
  wire [5:0] _foundTLB_T_1814 = _foundTLB_T_1813 | _foundTLB_T_1783;
  wire [5:0] _foundTLB_T_1784 = tlbHit_20_1 ? tlb_20_PS : 6'h0;
  wire [5:0] _foundTLB_T_1815 = _foundTLB_T_1814 | _foundTLB_T_1784;
  wire [5:0] _foundTLB_T_1785 = tlbHit_21_1 ? tlb_21_PS : 6'h0;
  wire [5:0] _foundTLB_T_1816 = _foundTLB_T_1815 | _foundTLB_T_1785;
  wire [5:0] _foundTLB_T_1786 = tlbHit_22_1 ? tlb_22_PS : 6'h0;
  wire [5:0] _foundTLB_T_1817 = _foundTLB_T_1816 | _foundTLB_T_1786;
  wire [5:0] _foundTLB_T_1787 = tlbHit_23_1 ? tlb_23_PS : 6'h0;
  wire [5:0] _foundTLB_T_1818 = _foundTLB_T_1817 | _foundTLB_T_1787;
  wire [5:0] _foundTLB_T_1788 = tlbHit_24_1 ? tlb_24_PS : 6'h0;
  wire [5:0] _foundTLB_T_1819 = _foundTLB_T_1818 | _foundTLB_T_1788;
  wire [5:0] _foundTLB_T_1789 = tlbHit_25_1 ? tlb_25_PS : 6'h0;
  wire [5:0] _foundTLB_T_1820 = _foundTLB_T_1819 | _foundTLB_T_1789;
  wire [5:0] _foundTLB_T_1790 = tlbHit_26_1 ? tlb_26_PS : 6'h0;
  wire [5:0] _foundTLB_T_1821 = _foundTLB_T_1820 | _foundTLB_T_1790;
  wire [5:0] _foundTLB_T_1791 = tlbHit_27_1 ? tlb_27_PS : 6'h0;
  wire [5:0] _foundTLB_T_1822 = _foundTLB_T_1821 | _foundTLB_T_1791;
  wire [5:0] _foundTLB_T_1792 = tlbHit_28_1 ? tlb_28_PS : 6'h0;
  wire [5:0] _foundTLB_T_1823 = _foundTLB_T_1822 | _foundTLB_T_1792;
  wire [5:0] _foundTLB_T_1793 = tlbHit_29_1 ? tlb_29_PS : 6'h0;
  wire [5:0] _foundTLB_T_1824 = _foundTLB_T_1823 | _foundTLB_T_1793;
  wire [5:0] _foundTLB_T_1794 = tlbHit_30_1 ? tlb_30_PS : 6'h0;
  wire [5:0] _foundTLB_T_1825 = _foundTLB_T_1824 | _foundTLB_T_1794;
  wire [5:0] _foundTLB_T_1795 = tlbHit_31_1 ? tlb_31_PS : 6'h0;
  wire [5:0] foundTLB_1_PS = _foundTLB_T_1825 | _foundTLB_T_1795;
  wire  _oddPG_T_3 = foundTLB_1_PS == 6'hc;
  wire  oddPG_1 = foundTLB_1_PS == 6'hc ? EXVA[12] : EXVA[22];
  wire  _foundTLB_T_960 = tlbHit_15_1 & tlb_15_P1_V;
  wire  _foundTLB_T_991 = tlbHit_0_1 & tlb_0_P1_V | tlbHit_1_1 & tlb_1_P1_V | tlbHit_2_1 & tlb_2_P1_V | tlbHit_3_1 &
    tlb_3_P1_V | tlbHit_4_1 & tlb_4_P1_V | tlbHit_5_1 & tlb_5_P1_V | tlbHit_6_1 & tlb_6_P1_V | tlbHit_7_1 & tlb_7_P1_V
     | tlbHit_8_1 & tlb_8_P1_V | tlbHit_9_1 & tlb_9_P1_V | tlbHit_10_1 & tlb_10_P1_V | tlbHit_11_1 & tlb_11_P1_V |
    tlbHit_12_1 & tlb_12_P1_V | tlbHit_13_1 & tlb_13_P1_V | tlbHit_14_1 & tlb_14_P1_V | _foundTLB_T_960;
  wire  _foundTLB_T_1006 = _foundTLB_T_991 | tlbHit_16_1 & tlb_16_P1_V | tlbHit_17_1 & tlb_17_P1_V | tlbHit_18_1 &
    tlb_18_P1_V | tlbHit_19_1 & tlb_19_P1_V | tlbHit_20_1 & tlb_20_P1_V | tlbHit_21_1 & tlb_21_P1_V | tlbHit_22_1 &
    tlb_22_P1_V | tlbHit_23_1 & tlb_23_P1_V | tlbHit_24_1 & tlb_24_P1_V | tlbHit_25_1 & tlb_25_P1_V | tlbHit_26_1 &
    tlb_26_P1_V | tlbHit_27_1 & tlb_27_P1_V | tlbHit_28_1 & tlb_28_P1_V | tlbHit_29_1 & tlb_29_P1_V | tlbHit_30_1 &
    tlb_30_P1_V;
  wire  foundTLB_1_P1_V = _foundTLB_T_1006 | tlbHit_31_1 & tlb_31_P1_V;
  wire  _foundTLB_T_1275 = tlbHit_15_1 & tlb_15_P0_V;
  wire  _foundTLB_T_1306 = tlbHit_0_1 & tlb_0_P0_V | tlbHit_1_1 & tlb_1_P0_V | tlbHit_2_1 & tlb_2_P0_V | tlbHit_3_1 &
    tlb_3_P0_V | tlbHit_4_1 & tlb_4_P0_V | tlbHit_5_1 & tlb_5_P0_V | tlbHit_6_1 & tlb_6_P0_V | tlbHit_7_1 & tlb_7_P0_V
     | tlbHit_8_1 & tlb_8_P0_V | tlbHit_9_1 & tlb_9_P0_V | tlbHit_10_1 & tlb_10_P0_V | tlbHit_11_1 & tlb_11_P0_V |
    tlbHit_12_1 & tlb_12_P0_V | tlbHit_13_1 & tlb_13_P0_V | tlbHit_14_1 & tlb_14_P0_V | _foundTLB_T_1275;
  wire  _foundTLB_T_1321 = _foundTLB_T_1306 | tlbHit_16_1 & tlb_16_P0_V | tlbHit_17_1 & tlb_17_P0_V | tlbHit_18_1 &
    tlb_18_P0_V | tlbHit_19_1 & tlb_19_P0_V | tlbHit_20_1 & tlb_20_P0_V | tlbHit_21_1 & tlb_21_P0_V | tlbHit_22_1 &
    tlb_22_P0_V | tlbHit_23_1 & tlb_23_P0_V | tlbHit_24_1 & tlb_24_P0_V | tlbHit_25_1 & tlb_25_P0_V | tlbHit_26_1 &
    tlb_26_P0_V | tlbHit_27_1 & tlb_27_P0_V | tlbHit_28_1 & tlb_28_P0_V | tlbHit_29_1 & tlb_29_P0_V | tlbHit_30_1 &
    tlb_30_P0_V;
  wire  foundTLB_1_P0_V = _foundTLB_T_1321 | tlbHit_31_1 & tlb_31_P0_V;
  wire  foundP_1_V = oddPG_1 ? foundTLB_1_P1_V : foundTLB_1_P0_V;
  wire  _GEN_71 = EXVA[31:29] == csrs_28_VSEG & (csrs_28_PLV0 & _T_11 | csrs_28_PLV3 & _T_13) ? 1'h0 : ~foundP_1_V;
  wire  invalid_1 = EXVA[31:29] == csrs_27_VSEG & (csrs_27_PLV0 & crmd_PLV == 2'h0 | csrs_27_PLV3 & crmd_PLV == 2'h3) ? 1'h0
     : _GEN_71;
  wire [1:0] _foundTLB_T_1134 = tlbHit_0_1 ? tlb_0_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1135 = tlbHit_1_1 ? tlb_1_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1166 = _foundTLB_T_1134 | _foundTLB_T_1135;
  wire [1:0] _foundTLB_T_1136 = tlbHit_2_1 ? tlb_2_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1167 = _foundTLB_T_1166 | _foundTLB_T_1136;
  wire [1:0] _foundTLB_T_1137 = tlbHit_3_1 ? tlb_3_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1168 = _foundTLB_T_1167 | _foundTLB_T_1137;
  wire [1:0] _foundTLB_T_1138 = tlbHit_4_1 ? tlb_4_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1169 = _foundTLB_T_1168 | _foundTLB_T_1138;
  wire [1:0] _foundTLB_T_1139 = tlbHit_5_1 ? tlb_5_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1170 = _foundTLB_T_1169 | _foundTLB_T_1139;
  wire [1:0] _foundTLB_T_1140 = tlbHit_6_1 ? tlb_6_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1171 = _foundTLB_T_1170 | _foundTLB_T_1140;
  wire [1:0] _foundTLB_T_1141 = tlbHit_7_1 ? tlb_7_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1172 = _foundTLB_T_1171 | _foundTLB_T_1141;
  wire [1:0] _foundTLB_T_1142 = tlbHit_8_1 ? tlb_8_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1173 = _foundTLB_T_1172 | _foundTLB_T_1142;
  wire [1:0] _foundTLB_T_1143 = tlbHit_9_1 ? tlb_9_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1174 = _foundTLB_T_1173 | _foundTLB_T_1143;
  wire [1:0] _foundTLB_T_1144 = tlbHit_10_1 ? tlb_10_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1175 = _foundTLB_T_1174 | _foundTLB_T_1144;
  wire [1:0] _foundTLB_T_1145 = tlbHit_11_1 ? tlb_11_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1176 = _foundTLB_T_1175 | _foundTLB_T_1145;
  wire [1:0] _foundTLB_T_1146 = tlbHit_12_1 ? tlb_12_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1177 = _foundTLB_T_1176 | _foundTLB_T_1146;
  wire [1:0] _foundTLB_T_1147 = tlbHit_13_1 ? tlb_13_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1178 = _foundTLB_T_1177 | _foundTLB_T_1147;
  wire [1:0] _foundTLB_T_1148 = tlbHit_14_1 ? tlb_14_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1179 = _foundTLB_T_1178 | _foundTLB_T_1148;
  wire [1:0] _foundTLB_T_1149 = tlbHit_15_1 ? tlb_15_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1180 = _foundTLB_T_1179 | _foundTLB_T_1149;
  wire [1:0] _foundTLB_T_1150 = tlbHit_16_1 ? tlb_16_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1181 = _foundTLB_T_1180 | _foundTLB_T_1150;
  wire [1:0] _foundTLB_T_1151 = tlbHit_17_1 ? tlb_17_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1182 = _foundTLB_T_1181 | _foundTLB_T_1151;
  wire [1:0] _foundTLB_T_1152 = tlbHit_18_1 ? tlb_18_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1183 = _foundTLB_T_1182 | _foundTLB_T_1152;
  wire [1:0] _foundTLB_T_1153 = tlbHit_19_1 ? tlb_19_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1184 = _foundTLB_T_1183 | _foundTLB_T_1153;
  wire [1:0] _foundTLB_T_1154 = tlbHit_20_1 ? tlb_20_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1185 = _foundTLB_T_1184 | _foundTLB_T_1154;
  wire [1:0] _foundTLB_T_1155 = tlbHit_21_1 ? tlb_21_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1186 = _foundTLB_T_1185 | _foundTLB_T_1155;
  wire [1:0] _foundTLB_T_1156 = tlbHit_22_1 ? tlb_22_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1187 = _foundTLB_T_1186 | _foundTLB_T_1156;
  wire [1:0] _foundTLB_T_1157 = tlbHit_23_1 ? tlb_23_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1188 = _foundTLB_T_1187 | _foundTLB_T_1157;
  wire [1:0] _foundTLB_T_1158 = tlbHit_24_1 ? tlb_24_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1189 = _foundTLB_T_1188 | _foundTLB_T_1158;
  wire [1:0] _foundTLB_T_1159 = tlbHit_25_1 ? tlb_25_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1190 = _foundTLB_T_1189 | _foundTLB_T_1159;
  wire [1:0] _foundTLB_T_1160 = tlbHit_26_1 ? tlb_26_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1191 = _foundTLB_T_1190 | _foundTLB_T_1160;
  wire [1:0] _foundTLB_T_1161 = tlbHit_27_1 ? tlb_27_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1192 = _foundTLB_T_1191 | _foundTLB_T_1161;
  wire [1:0] _foundTLB_T_1162 = tlbHit_28_1 ? tlb_28_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1193 = _foundTLB_T_1192 | _foundTLB_T_1162;
  wire [1:0] _foundTLB_T_1163 = tlbHit_29_1 ? tlb_29_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1194 = _foundTLB_T_1193 | _foundTLB_T_1163;
  wire [1:0] _foundTLB_T_1164 = tlbHit_30_1 ? tlb_30_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1195 = _foundTLB_T_1194 | _foundTLB_T_1164;
  wire [1:0] _foundTLB_T_1165 = tlbHit_31_1 ? tlb_31_P1_PLV : 2'h0;
  wire [1:0] foundTLB_1_P1_PLV = _foundTLB_T_1195 | _foundTLB_T_1165;
  wire [1:0] _foundTLB_T_1449 = tlbHit_0_1 ? tlb_0_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1450 = tlbHit_1_1 ? tlb_1_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1481 = _foundTLB_T_1449 | _foundTLB_T_1450;
  wire [1:0] _foundTLB_T_1451 = tlbHit_2_1 ? tlb_2_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1482 = _foundTLB_T_1481 | _foundTLB_T_1451;
  wire [1:0] _foundTLB_T_1452 = tlbHit_3_1 ? tlb_3_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1483 = _foundTLB_T_1482 | _foundTLB_T_1452;
  wire [1:0] _foundTLB_T_1453 = tlbHit_4_1 ? tlb_4_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1484 = _foundTLB_T_1483 | _foundTLB_T_1453;
  wire [1:0] _foundTLB_T_1454 = tlbHit_5_1 ? tlb_5_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1485 = _foundTLB_T_1484 | _foundTLB_T_1454;
  wire [1:0] _foundTLB_T_1455 = tlbHit_6_1 ? tlb_6_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1486 = _foundTLB_T_1485 | _foundTLB_T_1455;
  wire [1:0] _foundTLB_T_1456 = tlbHit_7_1 ? tlb_7_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1487 = _foundTLB_T_1486 | _foundTLB_T_1456;
  wire [1:0] _foundTLB_T_1457 = tlbHit_8_1 ? tlb_8_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1488 = _foundTLB_T_1487 | _foundTLB_T_1457;
  wire [1:0] _foundTLB_T_1458 = tlbHit_9_1 ? tlb_9_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1489 = _foundTLB_T_1488 | _foundTLB_T_1458;
  wire [1:0] _foundTLB_T_1459 = tlbHit_10_1 ? tlb_10_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1490 = _foundTLB_T_1489 | _foundTLB_T_1459;
  wire [1:0] _foundTLB_T_1460 = tlbHit_11_1 ? tlb_11_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1491 = _foundTLB_T_1490 | _foundTLB_T_1460;
  wire [1:0] _foundTLB_T_1461 = tlbHit_12_1 ? tlb_12_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1492 = _foundTLB_T_1491 | _foundTLB_T_1461;
  wire [1:0] _foundTLB_T_1462 = tlbHit_13_1 ? tlb_13_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1493 = _foundTLB_T_1492 | _foundTLB_T_1462;
  wire [1:0] _foundTLB_T_1463 = tlbHit_14_1 ? tlb_14_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1494 = _foundTLB_T_1493 | _foundTLB_T_1463;
  wire [1:0] _foundTLB_T_1464 = tlbHit_15_1 ? tlb_15_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1495 = _foundTLB_T_1494 | _foundTLB_T_1464;
  wire [1:0] _foundTLB_T_1465 = tlbHit_16_1 ? tlb_16_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1496 = _foundTLB_T_1495 | _foundTLB_T_1465;
  wire [1:0] _foundTLB_T_1466 = tlbHit_17_1 ? tlb_17_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1497 = _foundTLB_T_1496 | _foundTLB_T_1466;
  wire [1:0] _foundTLB_T_1467 = tlbHit_18_1 ? tlb_18_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1498 = _foundTLB_T_1497 | _foundTLB_T_1467;
  wire [1:0] _foundTLB_T_1468 = tlbHit_19_1 ? tlb_19_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1499 = _foundTLB_T_1498 | _foundTLB_T_1468;
  wire [1:0] _foundTLB_T_1469 = tlbHit_20_1 ? tlb_20_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1500 = _foundTLB_T_1499 | _foundTLB_T_1469;
  wire [1:0] _foundTLB_T_1470 = tlbHit_21_1 ? tlb_21_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1501 = _foundTLB_T_1500 | _foundTLB_T_1470;
  wire [1:0] _foundTLB_T_1471 = tlbHit_22_1 ? tlb_22_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1502 = _foundTLB_T_1501 | _foundTLB_T_1471;
  wire [1:0] _foundTLB_T_1472 = tlbHit_23_1 ? tlb_23_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1503 = _foundTLB_T_1502 | _foundTLB_T_1472;
  wire [1:0] _foundTLB_T_1473 = tlbHit_24_1 ? tlb_24_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1504 = _foundTLB_T_1503 | _foundTLB_T_1473;
  wire [1:0] _foundTLB_T_1474 = tlbHit_25_1 ? tlb_25_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1505 = _foundTLB_T_1504 | _foundTLB_T_1474;
  wire [1:0] _foundTLB_T_1475 = tlbHit_26_1 ? tlb_26_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1506 = _foundTLB_T_1505 | _foundTLB_T_1475;
  wire [1:0] _foundTLB_T_1476 = tlbHit_27_1 ? tlb_27_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1507 = _foundTLB_T_1506 | _foundTLB_T_1476;
  wire [1:0] _foundTLB_T_1477 = tlbHit_28_1 ? tlb_28_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1508 = _foundTLB_T_1507 | _foundTLB_T_1477;
  wire [1:0] _foundTLB_T_1478 = tlbHit_29_1 ? tlb_29_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1509 = _foundTLB_T_1508 | _foundTLB_T_1478;
  wire [1:0] _foundTLB_T_1479 = tlbHit_30_1 ? tlb_30_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_1510 = _foundTLB_T_1509 | _foundTLB_T_1479;
  wire [1:0] _foundTLB_T_1480 = tlbHit_31_1 ? tlb_31_P0_PLV : 2'h0;
  wire [1:0] foundTLB_1_P0_PLV = _foundTLB_T_1510 | _foundTLB_T_1480;
  wire [1:0] foundP_1_PLV = oddPG_1 ? foundTLB_1_P1_PLV : foundTLB_1_P0_PLV;
  wire  _GEN_72 = EXVA[31:29] == csrs_28_VSEG & (csrs_28_PLV0 & _T_11 | csrs_28_PLV3 & _T_13) ? 1'h0 : crmd_PLV >
    foundP_1_PLV;
  wire  ppi_1 = EXVA[31:29] == csrs_27_VSEG & (csrs_27_PLV0 & crmd_PLV == 2'h0 | csrs_27_PLV3 & crmd_PLV == 2'h3) ? 1'h0
     : _GEN_72;
  reg  tlb_0_P1_D;
  reg  tlb_1_P1_D;
  reg  tlb_2_P1_D;
  reg  tlb_3_P1_D;
  reg  tlb_4_P1_D;
  reg  tlb_5_P1_D;
  reg  tlb_6_P1_D;
  reg  tlb_7_P1_D;
  reg  tlb_8_P1_D;
  reg  tlb_9_P1_D;
  reg  tlb_10_P1_D;
  reg  tlb_11_P1_D;
  reg  tlb_12_P1_D;
  reg  tlb_13_P1_D;
  reg  tlb_14_P1_D;
  reg  tlb_15_P1_D;
  wire  _foundTLB_T_1023 = tlbHit_15_1 & tlb_15_P1_D;
  wire  _foundTLB_T_1054 = tlbHit_0_1 & tlb_0_P1_D | tlbHit_1_1 & tlb_1_P1_D | tlbHit_2_1 & tlb_2_P1_D | tlbHit_3_1 &
    tlb_3_P1_D | tlbHit_4_1 & tlb_4_P1_D | tlbHit_5_1 & tlb_5_P1_D | tlbHit_6_1 & tlb_6_P1_D | tlbHit_7_1 & tlb_7_P1_D
     | tlbHit_8_1 & tlb_8_P1_D | tlbHit_9_1 & tlb_9_P1_D | tlbHit_10_1 & tlb_10_P1_D | tlbHit_11_1 & tlb_11_P1_D |
    tlbHit_12_1 & tlb_12_P1_D | tlbHit_13_1 & tlb_13_P1_D | tlbHit_14_1 & tlb_14_P1_D | _foundTLB_T_1023;
  reg  tlb_16_P1_D;
  reg  tlb_17_P1_D;
  reg  tlb_18_P1_D;
  reg  tlb_19_P1_D;
  reg  tlb_20_P1_D;
  reg  tlb_21_P1_D;
  reg  tlb_22_P1_D;
  reg  tlb_23_P1_D;
  reg  tlb_24_P1_D;
  reg  tlb_25_P1_D;
  reg  tlb_26_P1_D;
  reg  tlb_27_P1_D;
  reg  tlb_28_P1_D;
  reg  tlb_29_P1_D;
  reg  tlb_30_P1_D;
  wire  _foundTLB_T_1069 = _foundTLB_T_1054 | tlbHit_16_1 & tlb_16_P1_D | tlbHit_17_1 & tlb_17_P1_D | tlbHit_18_1 &
    tlb_18_P1_D | tlbHit_19_1 & tlb_19_P1_D | tlbHit_20_1 & tlb_20_P1_D | tlbHit_21_1 & tlb_21_P1_D | tlbHit_22_1 &
    tlb_22_P1_D | tlbHit_23_1 & tlb_23_P1_D | tlbHit_24_1 & tlb_24_P1_D | tlbHit_25_1 & tlb_25_P1_D | tlbHit_26_1 &
    tlb_26_P1_D | tlbHit_27_1 & tlb_27_P1_D | tlbHit_28_1 & tlb_28_P1_D | tlbHit_29_1 & tlb_29_P1_D | tlbHit_30_1 &
    tlb_30_P1_D;
  reg  tlb_31_P1_D;
  wire  foundTLB_1_P1_D = _foundTLB_T_1069 | tlbHit_31_1 & tlb_31_P1_D;
  reg  tlb_0_P0_D;
  reg  tlb_1_P0_D;
  reg  tlb_2_P0_D;
  reg  tlb_3_P0_D;
  reg  tlb_4_P0_D;
  reg  tlb_5_P0_D;
  reg  tlb_6_P0_D;
  reg  tlb_7_P0_D;
  reg  tlb_8_P0_D;
  reg  tlb_9_P0_D;
  reg  tlb_10_P0_D;
  reg  tlb_11_P0_D;
  reg  tlb_12_P0_D;
  reg  tlb_13_P0_D;
  reg  tlb_14_P0_D;
  reg  tlb_15_P0_D;
  wire  _foundTLB_T_1338 = tlbHit_15_1 & tlb_15_P0_D;
  wire  _foundTLB_T_1369 = tlbHit_0_1 & tlb_0_P0_D | tlbHit_1_1 & tlb_1_P0_D | tlbHit_2_1 & tlb_2_P0_D | tlbHit_3_1 &
    tlb_3_P0_D | tlbHit_4_1 & tlb_4_P0_D | tlbHit_5_1 & tlb_5_P0_D | tlbHit_6_1 & tlb_6_P0_D | tlbHit_7_1 & tlb_7_P0_D
     | tlbHit_8_1 & tlb_8_P0_D | tlbHit_9_1 & tlb_9_P0_D | tlbHit_10_1 & tlb_10_P0_D | tlbHit_11_1 & tlb_11_P0_D |
    tlbHit_12_1 & tlb_12_P0_D | tlbHit_13_1 & tlb_13_P0_D | tlbHit_14_1 & tlb_14_P0_D | _foundTLB_T_1338;
  reg  tlb_16_P0_D;
  reg  tlb_17_P0_D;
  reg  tlb_18_P0_D;
  reg  tlb_19_P0_D;
  reg  tlb_20_P0_D;
  reg  tlb_21_P0_D;
  reg  tlb_22_P0_D;
  reg  tlb_23_P0_D;
  reg  tlb_24_P0_D;
  reg  tlb_25_P0_D;
  reg  tlb_26_P0_D;
  reg  tlb_27_P0_D;
  reg  tlb_28_P0_D;
  reg  tlb_29_P0_D;
  reg  tlb_30_P0_D;
  wire  _foundTLB_T_1384 = _foundTLB_T_1369 | tlbHit_16_1 & tlb_16_P0_D | tlbHit_17_1 & tlb_17_P0_D | tlbHit_18_1 &
    tlb_18_P0_D | tlbHit_19_1 & tlb_19_P0_D | tlbHit_20_1 & tlb_20_P0_D | tlbHit_21_1 & tlb_21_P0_D | tlbHit_22_1 &
    tlb_22_P0_D | tlbHit_23_1 & tlb_23_P0_D | tlbHit_24_1 & tlb_24_P0_D | tlbHit_25_1 & tlb_25_P0_D | tlbHit_26_1 &
    tlb_26_P0_D | tlbHit_27_1 & tlb_27_P0_D | tlbHit_28_1 & tlb_28_P0_D | tlbHit_29_1 & tlb_29_P0_D | tlbHit_30_1 &
    tlb_30_P0_D;
  reg  tlb_31_P0_D;
  wire  foundTLB_1_P0_D = _foundTLB_T_1384 | tlbHit_31_1 & tlb_31_P0_D;
  wire  foundP_1_D = oddPG_1 ? foundTLB_1_P1_D : foundTLB_1_P0_D;
  wire  _GEN_73 = EXVA[31:29] == csrs_28_VSEG & (csrs_28_PLV0 & _T_11 | csrs_28_PLV3 & _T_13) ? 1'h0 : ~foundP_1_D;
  wire  pme_1 = EXVA[31:29] == csrs_27_VSEG & (csrs_27_PLV0 & crmd_PLV == 2'h0 | csrs_27_PLV3 & crmd_PLV == 2'h3) ? 1'h0
     : _GEN_73;
  wire [1:0] _T_629 = _T_138 ? 2'h1 : 2'h0;
  wire [1:0] _T_630 = _T_136 ? 2'h1 : _T_629;
  wire [1:0] _T_631 = _T_134 ? 2'h1 : _T_630;
  wire [1:0] _T_632 = _T_132 ? 2'h0 : _T_631;
  wire [1:0] _T_633 = _T_130 ? 2'h0 : _T_632;
  wire [1:0] _T_634 = _T_128 ? 2'h0 : _T_633;
  wire [1:0] _T_635 = _T_126 ? 2'h3 : _T_634;
  wire [1:0] _T_636 = _T_124 ? 2'h2 : _T_635;
  wire [1:0] _T_637 = _T_122 ? 2'h0 : _T_636;
  wire [1:0] _T_638 = _T_120 ? 2'h0 : _T_637;
  wire [1:0] _T_639 = _T_118 ? 2'h0 : _T_638;
  wire [1:0] _T_640 = _T_116 ? 2'h0 : _T_639;
  wire [1:0] _T_641 = _T_114 ? 2'h0 : _T_640;
  wire [1:0] _T_642 = _T_112 ? 2'h0 : _T_641;
  wire [1:0] _T_643 = _T_110 ? 2'h0 : _T_642;
  wire [1:0] _T_644 = _T_108 ? 2'h0 : _T_643;
  wire [1:0] _T_645 = _T_106 ? 2'h0 : _T_644;
  wire [1:0] _T_646 = _T_104 ? 2'h0 : _T_645;
  wire [1:0] _T_647 = _T_102 ? 2'h0 : _T_646;
  wire [1:0] _T_648 = _T_100 ? 2'h0 : _T_647;
  wire [1:0] _T_649 = _T_98 ? 2'h0 : _T_648;
  wire [1:0] _T_650 = _T_96 ? 2'h0 : _T_649;
  wire [1:0] _T_651 = _T_94 ? 2'h0 : _T_650;
  wire [1:0] _T_652 = _T_92 ? 2'h0 : _T_651;
  wire [1:0] _T_653 = _T_90 ? 2'h0 : _T_652;
  wire [1:0] _T_654 = _T_88 ? 2'h0 : _T_653;
  wire [1:0] _T_655 = _T_86 ? 2'h0 : _T_654;
  wire [1:0] _T_656 = _T_84 ? 2'h0 : _T_655;
  wire [1:0] _T_657 = _T_82 ? 2'h0 : _T_656;
  wire [1:0] _T_658 = _T_80 ? 2'h0 : _T_657;
  wire [1:0] _T_659 = _T_78 ? 2'h0 : _T_658;
  wire [1:0] _T_660 = _T_76 ? 2'h0 : _T_659;
  wire [1:0] _T_661 = _T_74 ? 2'h0 : _T_660;
  wire [1:0] _T_662 = _T_72 ? 2'h0 : _T_661;
  wire [1:0] _T_663 = _T_70 ? 2'h0 : _T_662;
  wire [1:0] _T_664 = _T_68 ? 2'h0 : _T_663;
  wire [1:0] _T_665 = _T_66 ? 2'h0 : _T_664;
  wire [1:0] _T_666 = _T_64 ? 2'h0 : _T_665;
  wire [1:0] _T_667 = _T_62 ? 2'h0 : _T_666;
  wire [1:0] _T_668 = _T_60 ? 2'h0 : _T_667;
  wire [1:0] _T_669 = _T_58 ? 2'h0 : _T_668;
  wire [1:0] _T_670 = _T_56 ? 2'h0 : _T_669;
  wire [1:0] _T_671 = _T_54 ? 2'h0 : _T_670;
  wire [1:0] _T_672 = _T_52 ? 2'h0 : _T_671;
  wire [1:0] _T_673 = _T_50 ? 2'h0 : _T_672;
  wire [1:0] _T_674 = _T_48 ? 2'h0 : _T_673;
  wire [1:0] _T_675 = _T_46 ? 2'h0 : _T_674;
  wire [1:0] _T_676 = _T_44 ? 2'h0 : _T_675;
  wire [1:0] _T_677 = _T_42 ? 2'h0 : _T_676;
  wire [1:0] _T_678 = _T_40 ? 2'h0 : _T_677;
  wire [1:0] c0_2 = _T_38 ? 2'h0 : _T_678;
  wire  _GEN_87 = pme_1 & c0_2[0] & _lo_T_2;
  wire  _GEN_91 = ppi_1 ? 1'h0 : _GEN_87;
  wire  _GEN_97 = invalid_1 ? 1'h0 : _GEN_91;
  wire  _GEN_104 = miss_1 ? 1'h0 : _GEN_97;
  wire  _GEN_112 = crmd_DA ? 1'h0 : _GEN_104;
  wire  _GEN_120 = memADEM ? 1'h0 : _GEN_112;
  wire  _GEN_129 = memALE ? 1'h0 : _GEN_120;
  wire  _GEN_138 = c0_3 == 3'h7 | c0_11 & d[4:3] != 2'h2 ? 1'h0 : _GEN_129;
  wire  _GEN_152 = ID_OK & _GEN_138;
  wire  PME = dStallReg ? 1'h0 : _GEN_152;
  wire  _GEN_23 = invalid ? 1'h0 : ppi;
  wire  _GEN_27 = miss ? 1'h0 : _GEN_23;
  wire  _GEN_32 = crmd_DA ? 1'h0 : _GEN_27;
  wire  _GEN_37 = PC[1:0] != 2'h0 | PC[31] & crmd_PLV != 2'h0 ? 1'h0 : _GEN_32;
  wire  _GEN_42 = ~INT & ~idle & _GEN_37;
  wire  _GEN_47 = dStallReg | iStallReg ? 1'h0 : _GEN_42;
  wire  _GEN_90 = ppi_1 ? _lo_T_2 : _GEN_47;
  wire  _GEN_96 = invalid_1 ? _GEN_47 : _GEN_90;
  wire  _GEN_103 = miss_1 ? _GEN_47 : _GEN_96;
  wire  _GEN_111 = crmd_DA ? _GEN_47 : _GEN_103;
  wire  _GEN_119 = memADEM ? _GEN_47 : _GEN_111;
  wire  _GEN_128 = memALE ? _GEN_47 : _GEN_119;
  wire  _GEN_137 = c0_3 == 3'h7 | c0_11 & d[4:3] != 2'h2 ? _GEN_47 : _GEN_128;
  wire  _GEN_151 = ID_OK ? _GEN_137 : _GEN_47;
  wire  PPI = dStallReg ? _GEN_47 : _GEN_151;
  wire  _GEN_85 = c0_2[0] & _lo_T_2;
  wire  _GEN_94 = invalid_1 & _GEN_85;
  wire  _GEN_101 = miss_1 ? 1'h0 : _GEN_94;
  wire  _GEN_109 = crmd_DA ? 1'h0 : _GEN_101;
  wire  _GEN_117 = memADEM ? 1'h0 : _GEN_109;
  wire  _GEN_126 = memALE ? 1'h0 : _GEN_117;
  wire  _GEN_135 = c0_3 == 3'h7 | c0_11 & d[4:3] != 2'h2 ? 1'h0 : _GEN_126;
  wire  _GEN_149 = ID_OK & _GEN_135;
  wire  PIS = dStallReg ? 1'h0 : _GEN_149;
  wire  _GEN_26 = miss ? 1'h0 : invalid;
  wire  _GEN_31 = crmd_DA ? 1'h0 : _GEN_26;
  wire  _GEN_36 = PC[1:0] != 2'h0 | PC[31] & crmd_PLV != 2'h0 ? 1'h0 : _GEN_31;
  wire  _GEN_41 = ~INT & ~idle & _GEN_36;
  wire  PIF = dStallReg | iStallReg ? 1'h0 : _GEN_41;
  wire  _GEN_86 = c0_2[0] ? 1'h0 : _lo_T_2;
  wire  _GEN_95 = invalid_1 & _GEN_86;
  wire  _GEN_102 = miss_1 ? 1'h0 : _GEN_95;
  wire  _GEN_110 = crmd_DA ? 1'h0 : _GEN_102;
  wire  _GEN_118 = memADEM ? 1'h0 : _GEN_110;
  wire  _GEN_127 = memALE ? 1'h0 : _GEN_118;
  wire  _GEN_136 = c0_3 == 3'h7 | c0_11 & d[4:3] != 2'h2 ? 1'h0 : _GEN_127;
  wire  _GEN_150 = ID_OK & _GEN_136;
  wire  PIL = dStallReg ? 1'h0 : _GEN_150;
  wire [15:0] _excp_T = {INT,PIL,PIS,PIF,PME,PPI,ADEF,ADEM,excp_lo};
  wire  excp = |_excp_T;
  reg [19:0] tlb_0_P0_PPN;
  reg [1:0] tlb_0_P0_MAT;
  reg [19:0] tlb_0_P1_PPN;
  reg [1:0] tlb_0_P1_MAT;
  reg [19:0] tlb_1_P0_PPN;
  reg [1:0] tlb_1_P0_MAT;
  reg [19:0] tlb_1_P1_PPN;
  reg [1:0] tlb_1_P1_MAT;
  reg [19:0] tlb_2_P0_PPN;
  reg [1:0] tlb_2_P0_MAT;
  reg [19:0] tlb_2_P1_PPN;
  reg [1:0] tlb_2_P1_MAT;
  reg [19:0] tlb_3_P0_PPN;
  reg [1:0] tlb_3_P0_MAT;
  reg [19:0] tlb_3_P1_PPN;
  reg [1:0] tlb_3_P1_MAT;
  reg [19:0] tlb_4_P0_PPN;
  reg [1:0] tlb_4_P0_MAT;
  reg [19:0] tlb_4_P1_PPN;
  reg [1:0] tlb_4_P1_MAT;
  reg [19:0] tlb_5_P0_PPN;
  reg [1:0] tlb_5_P0_MAT;
  reg [19:0] tlb_5_P1_PPN;
  reg [1:0] tlb_5_P1_MAT;
  reg [19:0] tlb_6_P0_PPN;
  reg [1:0] tlb_6_P0_MAT;
  reg [19:0] tlb_6_P1_PPN;
  reg [1:0] tlb_6_P1_MAT;
  reg [19:0] tlb_7_P0_PPN;
  reg [1:0] tlb_7_P0_MAT;
  reg [19:0] tlb_7_P1_PPN;
  reg [1:0] tlb_7_P1_MAT;
  reg [19:0] tlb_8_P0_PPN;
  reg [1:0] tlb_8_P0_MAT;
  reg [19:0] tlb_8_P1_PPN;
  reg [1:0] tlb_8_P1_MAT;
  reg [19:0] tlb_9_P0_PPN;
  reg [1:0] tlb_9_P0_MAT;
  reg [19:0] tlb_9_P1_PPN;
  reg [1:0] tlb_9_P1_MAT;
  reg [19:0] tlb_10_P0_PPN;
  reg [1:0] tlb_10_P0_MAT;
  reg [19:0] tlb_10_P1_PPN;
  reg [1:0] tlb_10_P1_MAT;
  reg [19:0] tlb_11_P0_PPN;
  reg [1:0] tlb_11_P0_MAT;
  reg [19:0] tlb_11_P1_PPN;
  reg [1:0] tlb_11_P1_MAT;
  reg [19:0] tlb_12_P0_PPN;
  reg [1:0] tlb_12_P0_MAT;
  reg [19:0] tlb_12_P1_PPN;
  reg [1:0] tlb_12_P1_MAT;
  reg [19:0] tlb_13_P0_PPN;
  reg [1:0] tlb_13_P0_MAT;
  reg [19:0] tlb_13_P1_PPN;
  reg [1:0] tlb_13_P1_MAT;
  reg [19:0] tlb_14_P0_PPN;
  reg [1:0] tlb_14_P0_MAT;
  reg [19:0] tlb_14_P1_PPN;
  reg [1:0] tlb_14_P1_MAT;
  reg [19:0] tlb_15_P0_PPN;
  reg [1:0] tlb_15_P0_MAT;
  reg [19:0] tlb_15_P1_PPN;
  reg [1:0] tlb_15_P1_MAT;
  reg [19:0] tlb_16_P0_PPN;
  reg [1:0] tlb_16_P0_MAT;
  reg [19:0] tlb_16_P1_PPN;
  reg [1:0] tlb_16_P1_MAT;
  reg [19:0] tlb_17_P0_PPN;
  reg [1:0] tlb_17_P0_MAT;
  reg [19:0] tlb_17_P1_PPN;
  reg [1:0] tlb_17_P1_MAT;
  reg [19:0] tlb_18_P0_PPN;
  reg [1:0] tlb_18_P0_MAT;
  reg [19:0] tlb_18_P1_PPN;
  reg [1:0] tlb_18_P1_MAT;
  reg [19:0] tlb_19_P0_PPN;
  reg [1:0] tlb_19_P0_MAT;
  reg [19:0] tlb_19_P1_PPN;
  reg [1:0] tlb_19_P1_MAT;
  reg [19:0] tlb_20_P0_PPN;
  reg [1:0] tlb_20_P0_MAT;
  reg [19:0] tlb_20_P1_PPN;
  reg [1:0] tlb_20_P1_MAT;
  reg [19:0] tlb_21_P0_PPN;
  reg [1:0] tlb_21_P0_MAT;
  reg [19:0] tlb_21_P1_PPN;
  reg [1:0] tlb_21_P1_MAT;
  reg [19:0] tlb_22_P0_PPN;
  reg [1:0] tlb_22_P0_MAT;
  reg [19:0] tlb_22_P1_PPN;
  reg [1:0] tlb_22_P1_MAT;
  reg [19:0] tlb_23_P0_PPN;
  reg [1:0] tlb_23_P0_MAT;
  reg [19:0] tlb_23_P1_PPN;
  reg [1:0] tlb_23_P1_MAT;
  reg [19:0] tlb_24_P0_PPN;
  reg [1:0] tlb_24_P0_MAT;
  reg [19:0] tlb_24_P1_PPN;
  reg [1:0] tlb_24_P1_MAT;
  reg [19:0] tlb_25_P0_PPN;
  reg [1:0] tlb_25_P0_MAT;
  reg [19:0] tlb_25_P1_PPN;
  reg [1:0] tlb_25_P1_MAT;
  reg [19:0] tlb_26_P0_PPN;
  reg [1:0] tlb_26_P0_MAT;
  reg [19:0] tlb_26_P1_PPN;
  reg [1:0] tlb_26_P1_MAT;
  reg [19:0] tlb_27_P0_PPN;
  reg [1:0] tlb_27_P0_MAT;
  reg [19:0] tlb_27_P1_PPN;
  reg [1:0] tlb_27_P1_MAT;
  reg [19:0] tlb_28_P0_PPN;
  reg [1:0] tlb_28_P0_MAT;
  reg [19:0] tlb_28_P1_PPN;
  reg [1:0] tlb_28_P1_MAT;
  reg [19:0] tlb_29_P0_PPN;
  reg [1:0] tlb_29_P0_MAT;
  reg [19:0] tlb_29_P1_PPN;
  reg [1:0] tlb_29_P1_MAT;
  reg [19:0] tlb_30_P0_PPN;
  reg [1:0] tlb_30_P0_MAT;
  reg [19:0] tlb_30_P1_PPN;
  reg [1:0] tlb_30_P1_MAT;
  reg [19:0] tlb_31_P0_PPN;
  reg [1:0] tlb_31_P0_MAT;
  reg [19:0] tlb_31_P1_PPN;
  reg [1:0] tlb_31_P1_MAT;
  wire [28:0] pa_lo = PC[28:0];
  wire [31:0] _pa_T = {csrs_27_PSEG,pa_lo};
  wire [31:0] _pa_T_1 = {csrs_28_PSEG,pa_lo};
  wire [19:0] _foundTLB_T_252 = tlbHit_0 ? tlb_0_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_253 = tlbHit_1 ? tlb_1_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_254 = tlbHit_2 ? tlb_2_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_255 = tlbHit_3 ? tlb_3_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_256 = tlbHit_4 ? tlb_4_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_257 = tlbHit_5 ? tlb_5_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_258 = tlbHit_6 ? tlb_6_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_259 = tlbHit_7 ? tlb_7_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_260 = tlbHit_8 ? tlb_8_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_261 = tlbHit_9 ? tlb_9_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_262 = tlbHit_10 ? tlb_10_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_263 = tlbHit_11 ? tlb_11_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_264 = tlbHit_12 ? tlb_12_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_265 = tlbHit_13 ? tlb_13_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_266 = tlbHit_14 ? tlb_14_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_267 = tlbHit_15 ? tlb_15_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_268 = tlbHit_16 ? tlb_16_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_269 = tlbHit_17 ? tlb_17_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_270 = tlbHit_18 ? tlb_18_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_271 = tlbHit_19 ? tlb_19_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_272 = tlbHit_20 ? tlb_20_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_273 = tlbHit_21 ? tlb_21_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_274 = tlbHit_22 ? tlb_22_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_275 = tlbHit_23 ? tlb_23_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_276 = tlbHit_24 ? tlb_24_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_277 = tlbHit_25 ? tlb_25_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_278 = tlbHit_26 ? tlb_26_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_279 = tlbHit_27 ? tlb_27_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_280 = tlbHit_28 ? tlb_28_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_281 = tlbHit_29 ? tlb_29_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_282 = tlbHit_30 ? tlb_30_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_283 = tlbHit_31 ? tlb_31_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_284 = _foundTLB_T_252 | _foundTLB_T_253;
  wire [19:0] _foundTLB_T_285 = _foundTLB_T_284 | _foundTLB_T_254;
  wire [19:0] _foundTLB_T_286 = _foundTLB_T_285 | _foundTLB_T_255;
  wire [19:0] _foundTLB_T_287 = _foundTLB_T_286 | _foundTLB_T_256;
  wire [19:0] _foundTLB_T_288 = _foundTLB_T_287 | _foundTLB_T_257;
  wire [19:0] _foundTLB_T_289 = _foundTLB_T_288 | _foundTLB_T_258;
  wire [19:0] _foundTLB_T_290 = _foundTLB_T_289 | _foundTLB_T_259;
  wire [19:0] _foundTLB_T_291 = _foundTLB_T_290 | _foundTLB_T_260;
  wire [19:0] _foundTLB_T_292 = _foundTLB_T_291 | _foundTLB_T_261;
  wire [19:0] _foundTLB_T_293 = _foundTLB_T_292 | _foundTLB_T_262;
  wire [19:0] _foundTLB_T_294 = _foundTLB_T_293 | _foundTLB_T_263;
  wire [19:0] _foundTLB_T_295 = _foundTLB_T_294 | _foundTLB_T_264;
  wire [19:0] _foundTLB_T_296 = _foundTLB_T_295 | _foundTLB_T_265;
  wire [19:0] _foundTLB_T_297 = _foundTLB_T_296 | _foundTLB_T_266;
  wire [19:0] _foundTLB_T_298 = _foundTLB_T_297 | _foundTLB_T_267;
  wire [19:0] _foundTLB_T_299 = _foundTLB_T_298 | _foundTLB_T_268;
  wire [19:0] _foundTLB_T_300 = _foundTLB_T_299 | _foundTLB_T_269;
  wire [19:0] _foundTLB_T_301 = _foundTLB_T_300 | _foundTLB_T_270;
  wire [19:0] _foundTLB_T_302 = _foundTLB_T_301 | _foundTLB_T_271;
  wire [19:0] _foundTLB_T_303 = _foundTLB_T_302 | _foundTLB_T_272;
  wire [19:0] _foundTLB_T_304 = _foundTLB_T_303 | _foundTLB_T_273;
  wire [19:0] _foundTLB_T_305 = _foundTLB_T_304 | _foundTLB_T_274;
  wire [19:0] _foundTLB_T_306 = _foundTLB_T_305 | _foundTLB_T_275;
  wire [19:0] _foundTLB_T_307 = _foundTLB_T_306 | _foundTLB_T_276;
  wire [19:0] _foundTLB_T_308 = _foundTLB_T_307 | _foundTLB_T_277;
  wire [19:0] _foundTLB_T_309 = _foundTLB_T_308 | _foundTLB_T_278;
  wire [19:0] _foundTLB_T_310 = _foundTLB_T_309 | _foundTLB_T_279;
  wire [19:0] _foundTLB_T_311 = _foundTLB_T_310 | _foundTLB_T_280;
  wire [19:0] _foundTLB_T_312 = _foundTLB_T_311 | _foundTLB_T_281;
  wire [19:0] _foundTLB_T_313 = _foundTLB_T_312 | _foundTLB_T_282;
  wire [19:0] foundTLB_P1_PPN = _foundTLB_T_313 | _foundTLB_T_283;
  wire [19:0] _foundTLB_T_567 = tlbHit_0 ? tlb_0_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_568 = tlbHit_1 ? tlb_1_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_569 = tlbHit_2 ? tlb_2_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_570 = tlbHit_3 ? tlb_3_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_571 = tlbHit_4 ? tlb_4_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_572 = tlbHit_5 ? tlb_5_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_573 = tlbHit_6 ? tlb_6_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_574 = tlbHit_7 ? tlb_7_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_575 = tlbHit_8 ? tlb_8_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_576 = tlbHit_9 ? tlb_9_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_577 = tlbHit_10 ? tlb_10_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_578 = tlbHit_11 ? tlb_11_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_579 = tlbHit_12 ? tlb_12_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_580 = tlbHit_13 ? tlb_13_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_581 = tlbHit_14 ? tlb_14_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_582 = tlbHit_15 ? tlb_15_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_583 = tlbHit_16 ? tlb_16_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_584 = tlbHit_17 ? tlb_17_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_585 = tlbHit_18 ? tlb_18_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_586 = tlbHit_19 ? tlb_19_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_587 = tlbHit_20 ? tlb_20_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_588 = tlbHit_21 ? tlb_21_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_589 = tlbHit_22 ? tlb_22_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_590 = tlbHit_23 ? tlb_23_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_591 = tlbHit_24 ? tlb_24_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_592 = tlbHit_25 ? tlb_25_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_593 = tlbHit_26 ? tlb_26_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_594 = tlbHit_27 ? tlb_27_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_595 = tlbHit_28 ? tlb_28_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_596 = tlbHit_29 ? tlb_29_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_597 = tlbHit_30 ? tlb_30_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_598 = tlbHit_31 ? tlb_31_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_599 = _foundTLB_T_567 | _foundTLB_T_568;
  wire [19:0] _foundTLB_T_600 = _foundTLB_T_599 | _foundTLB_T_569;
  wire [19:0] _foundTLB_T_601 = _foundTLB_T_600 | _foundTLB_T_570;
  wire [19:0] _foundTLB_T_602 = _foundTLB_T_601 | _foundTLB_T_571;
  wire [19:0] _foundTLB_T_603 = _foundTLB_T_602 | _foundTLB_T_572;
  wire [19:0] _foundTLB_T_604 = _foundTLB_T_603 | _foundTLB_T_573;
  wire [19:0] _foundTLB_T_605 = _foundTLB_T_604 | _foundTLB_T_574;
  wire [19:0] _foundTLB_T_606 = _foundTLB_T_605 | _foundTLB_T_575;
  wire [19:0] _foundTLB_T_607 = _foundTLB_T_606 | _foundTLB_T_576;
  wire [19:0] _foundTLB_T_608 = _foundTLB_T_607 | _foundTLB_T_577;
  wire [19:0] _foundTLB_T_609 = _foundTLB_T_608 | _foundTLB_T_578;
  wire [19:0] _foundTLB_T_610 = _foundTLB_T_609 | _foundTLB_T_579;
  wire [19:0] _foundTLB_T_611 = _foundTLB_T_610 | _foundTLB_T_580;
  wire [19:0] _foundTLB_T_612 = _foundTLB_T_611 | _foundTLB_T_581;
  wire [19:0] _foundTLB_T_613 = _foundTLB_T_612 | _foundTLB_T_582;
  wire [19:0] _foundTLB_T_614 = _foundTLB_T_613 | _foundTLB_T_583;
  wire [19:0] _foundTLB_T_615 = _foundTLB_T_614 | _foundTLB_T_584;
  wire [19:0] _foundTLB_T_616 = _foundTLB_T_615 | _foundTLB_T_585;
  wire [19:0] _foundTLB_T_617 = _foundTLB_T_616 | _foundTLB_T_586;
  wire [19:0] _foundTLB_T_618 = _foundTLB_T_617 | _foundTLB_T_587;
  wire [19:0] _foundTLB_T_619 = _foundTLB_T_618 | _foundTLB_T_588;
  wire [19:0] _foundTLB_T_620 = _foundTLB_T_619 | _foundTLB_T_589;
  wire [19:0] _foundTLB_T_621 = _foundTLB_T_620 | _foundTLB_T_590;
  wire [19:0] _foundTLB_T_622 = _foundTLB_T_621 | _foundTLB_T_591;
  wire [19:0] _foundTLB_T_623 = _foundTLB_T_622 | _foundTLB_T_592;
  wire [19:0] _foundTLB_T_624 = _foundTLB_T_623 | _foundTLB_T_593;
  wire [19:0] _foundTLB_T_625 = _foundTLB_T_624 | _foundTLB_T_594;
  wire [19:0] _foundTLB_T_626 = _foundTLB_T_625 | _foundTLB_T_595;
  wire [19:0] _foundTLB_T_627 = _foundTLB_T_626 | _foundTLB_T_596;
  wire [19:0] _foundTLB_T_628 = _foundTLB_T_627 | _foundTLB_T_597;
  wire [19:0] foundTLB_P0_PPN = _foundTLB_T_628 | _foundTLB_T_598;
  wire [19:0] foundP_PPN = oddPG ? foundTLB_P1_PPN : foundTLB_P0_PPN;
  wire [11:0] pa_lo_2 = PC[11:0];
  wire [31:0] _pa_T_3 = {foundP_PPN,pa_lo_2};
  wire [9:0] pa_hi = foundP_PPN[19:10];
  wire [11:0] pa_lo_3 = PC[21:10];
  wire [21:0] _pa_T_4 = {pa_hi,pa_lo_3};
  wire [31:0] _pa_T_5 = _oddPG_T ? _pa_T_3 : {{10'd0}, _pa_T_4};
  wire [31:0] _GEN_8 = PC[31:29] == csrs_28_VSEG & (csrs_28_PLV0 & _T_11 | csrs_28_PLV3 & _T_13) ? _pa_T_1 : _pa_T_5;
  wire [31:0] pa = PC[31:29] == csrs_27_VSEG & (csrs_27_PLV0 & crmd_PLV == 2'h0 | csrs_27_PLV3 & crmd_PLV == 2'h3) ?
    _pa_T : _GEN_8;
  wire  _io_inst_req_valid_T_1 = ~dStallReg;
  wire [18:0] _GEN_48 = ~ADEF ? PC[31:13] : csrs_9_VPPN;
  wire [31:0] _GEN_49 = ~IF_OK ? PC : badv_VAddr;
  wire [18:0] _GEN_50 = ~IF_OK ? _GEN_48 : csrs_9_VPPN;
  wire [2:0] _T_493 = _T_154 ? 3'h2 : 3'h0;
  wire [2:0] _T_494 = _T_152 ? 3'h0 : _T_493;
  wire [2:0] _T_495 = _T_150 ? 3'h2 : _T_494;
  wire [2:0] _T_496 = _T_148 ? 3'h0 : _T_495;
  wire [2:0] _T_497 = _T_146 ? 3'h0 : _T_496;
  wire [2:0] _T_498 = _T_144 ? 3'h0 : _T_497;
  wire [2:0] _T_499 = _T_142 ? 3'h1 : _T_498;
  wire [2:0] _T_500 = _T_140 ? 3'h1 : _T_499;
  wire [2:0] _T_501 = _T_138 ? 3'h0 : _T_500;
  wire [2:0] _T_502 = _T_136 ? 3'h0 : _T_501;
  wire [2:0] _T_503 = _T_134 ? 3'h0 : _T_502;
  wire [2:0] _T_504 = _T_132 ? 3'h1 : _T_503;
  wire [2:0] _T_505 = _T_130 ? 3'h1 : _T_504;
  wire [2:0] _T_506 = _T_128 ? 3'h1 : _T_505;
  wire [2:0] _T_507 = _T_126 ? 3'h7 : _T_506;
  wire [2:0] _T_508 = _T_124 ? 3'h1 : _T_507;
  wire [2:0] _T_509 = _T_122 ? 3'h0 : _T_508;
  wire [2:0] _T_510 = _T_120 ? 3'h0 : _T_509;
  wire [2:0] _T_511 = _T_118 ? 3'h0 : _T_510;
  wire [2:0] _T_512 = _T_116 ? 3'h0 : _T_511;
  wire [2:0] _T_513 = _T_114 ? 3'h0 : _T_512;
  wire [2:0] _T_514 = _T_112 ? 3'h0 : _T_513;
  wire [2:0] _T_515 = _T_110 ? 3'h0 : _T_514;
  wire [2:0] _T_516 = _T_108 ? 3'h0 : _T_515;
  wire [2:0] _T_517 = _T_106 ? 3'h0 : _T_516;
  wire [2:0] _T_518 = _T_104 ? 3'h0 : _T_517;
  wire [2:0] _T_519 = _T_102 ? 3'h3 : _T_518;
  wire [2:0] _T_520 = _T_100 ? 3'h0 : _T_519;
  wire [2:0] _T_521 = _T_98 ? 3'h0 : _T_520;
  wire [2:0] _T_522 = _T_96 ? 3'h0 : _T_521;
  wire [2:0] _T_523 = _T_94 ? 3'h0 : _T_522;
  wire [2:0] _T_524 = _T_92 ? 3'h0 : _T_523;
  wire [2:0] _T_525 = _T_90 ? 3'h0 : _T_524;
  wire [2:0] _T_526 = _T_88 ? 3'h0 : _T_525;
  wire [2:0] _T_527 = _T_86 ? 3'h0 : _T_526;
  wire [2:0] _T_528 = _T_84 ? 3'h0 : _T_527;
  wire [2:0] _T_529 = _T_82 ? 3'h0 : _T_528;
  wire [2:0] _T_530 = _T_80 ? 3'h0 : _T_529;
  wire [2:0] _T_531 = _T_78 ? 3'h0 : _T_530;
  wire [2:0] _T_532 = _T_76 ? 3'h0 : _T_531;
  wire [2:0] _T_533 = _T_74 ? 3'h0 : _T_532;
  wire [2:0] _T_534 = _T_72 ? 3'h0 : _T_533;
  wire [2:0] _T_535 = _T_70 ? 3'h0 : _T_534;
  wire [2:0] _T_536 = _T_68 ? 3'h0 : _T_535;
  wire [2:0] _T_537 = _T_66 ? 3'h0 : _T_536;
  wire [2:0] _T_538 = _T_64 ? 3'h0 : _T_537;
  wire [2:0] _T_539 = _T_62 ? 3'h0 : _T_538;
  wire [2:0] _T_540 = _T_60 ? 3'h0 : _T_539;
  wire [2:0] _T_541 = _T_58 ? 3'h0 : _T_540;
  wire [2:0] _T_542 = _T_56 ? 3'h0 : _T_541;
  wire [2:0] _T_543 = _T_54 ? 3'h0 : _T_542;
  wire [2:0] _T_544 = _T_52 ? 3'h0 : _T_543;
  wire [2:0] _T_545 = _T_50 ? 3'h0 : _T_544;
  wire [2:0] _T_546 = _T_48 ? 3'h0 : _T_545;
  wire [2:0] _T_547 = _T_46 ? 3'h0 : _T_546;
  wire [2:0] _T_548 = _T_44 ? 3'h0 : _T_547;
  wire [2:0] _T_549 = _T_42 ? 3'h5 : _T_548;
  wire [2:0] _T_550 = _T_40 ? 3'h6 : _T_549;
  wire [2:0] c0_0 = _T_38 ? 3'h4 : _T_550;
  wire [1:0] _T_557 = _T_154 ? 2'h1 : 2'h0;
  wire [1:0] _T_558 = _T_152 ? 2'h0 : _T_557;
  wire [1:0] _T_559 = _T_150 ? 2'h2 : _T_558;
  wire [1:0] _T_560 = _T_148 ? 2'h0 : _T_559;
  wire [1:0] _T_561 = _T_146 ? 2'h0 : _T_560;
  wire [1:0] _T_562 = _T_144 ? 2'h0 : _T_561;
  wire [1:0] _T_563 = _T_142 ? 2'h2 : _T_562;
  wire [1:0] _T_564 = _T_140 ? 2'h2 : _T_563;
  wire [1:0] _T_565 = _T_138 ? 2'h0 : _T_564;
  wire [1:0] _T_566 = _T_136 ? 2'h0 : _T_565;
  wire [1:0] _T_567 = _T_134 ? 2'h0 : _T_566;
  wire [1:0] _T_568 = _T_132 ? 2'h2 : _T_567;
  wire [1:0] _T_569 = _T_130 ? 2'h2 : _T_568;
  wire [1:0] _T_570 = _T_128 ? 2'h2 : _T_569;
  wire [1:0] _T_571 = _T_126 ? 2'h2 : _T_570;
  wire [1:0] _T_572 = _T_124 ? 2'h2 : _T_571;
  wire [1:0] _T_573 = _T_122 ? 2'h2 : _T_572;
  wire [1:0] _T_574 = _T_120 ? 2'h2 : _T_573;
  wire [1:0] _T_575 = _T_118 ? 2'h0 : _T_574;
  wire [1:0] _T_576 = _T_116 ? 2'h0 : _T_575;
  wire [1:0] _T_577 = _T_114 ? 2'h0 : _T_576;
  wire [1:0] _T_578 = _T_112 ? 2'h0 : _T_577;
  wire [1:0] _T_579 = _T_110 ? 2'h0 : _T_578;
  wire [1:0] _T_580 = _T_108 ? 2'h0 : _T_579;
  wire [1:0] _T_581 = _T_106 ? 2'h0 : _T_580;
  wire [1:0] _T_582 = _T_104 ? 2'h0 : _T_581;
  wire [1:0] _T_583 = _T_102 ? 2'h2 : _T_582;
  wire [1:0] _T_584 = _T_100 ? 2'h2 : _T_583;
  wire [1:0] _T_585 = _T_98 ? 2'h2 : _T_584;
  wire [1:0] _T_586 = _T_96 ? 2'h2 : _T_585;
  wire [1:0] _T_587 = _T_94 ? 2'h2 : _T_586;
  wire [1:0] _T_588 = _T_92 ? 2'h2 : _T_587;
  wire [1:0] _T_589 = _T_90 ? 2'h2 : _T_588;
  wire [1:0] _T_590 = _T_88 ? 2'h2 : _T_589;
  wire [1:0] _T_591 = _T_86 ? 2'h2 : _T_590;
  wire [1:0] _T_592 = _T_84 ? 2'h2 : _T_591;
  wire [1:0] _T_593 = _T_82 ? 2'h0 : _T_592;
  wire [1:0] _T_594 = _T_80 ? 2'h0 : _T_593;
  wire [1:0] _T_595 = _T_78 ? 2'h2 : _T_594;
  wire [1:0] _T_596 = _T_76 ? 2'h2 : _T_595;
  wire [1:0] _T_597 = _T_74 ? 2'h2 : _T_596;
  wire [1:0] _T_598 = _T_72 ? 2'h2 : _T_597;
  wire [1:0] _T_599 = _T_70 ? 2'h2 : _T_598;
  wire [1:0] _T_600 = _T_68 ? 2'h2 : _T_599;
  wire [1:0] _T_601 = _T_66 ? 2'h2 : _T_600;
  wire [1:0] _T_602 = _T_64 ? 2'h2 : _T_601;
  wire [1:0] _T_603 = _T_62 ? 2'h2 : _T_602;
  wire [1:0] _T_604 = _T_60 ? 2'h2 : _T_603;
  wire [1:0] _T_605 = _T_58 ? 2'h2 : _T_604;
  wire [1:0] _T_606 = _T_56 ? 2'h2 : _T_605;
  wire [1:0] _T_607 = _T_54 ? 2'h2 : _T_606;
  wire [1:0] _T_608 = _T_52 ? 2'h2 : _T_607;
  wire [1:0] _T_609 = _T_50 ? 2'h2 : _T_608;
  wire [1:0] _T_610 = _T_48 ? 2'h2 : _T_609;
  wire [1:0] _T_611 = _T_46 ? 2'h2 : _T_610;
  wire [1:0] _T_612 = _T_44 ? 2'h2 : _T_611;
  wire [1:0] _T_613 = _T_42 ? 2'h2 : _T_612;
  wire [1:0] _T_614 = _T_40 ? 2'h2 : _T_613;
  wire [1:0] c0_1 = _T_38 ? 2'h3 : _T_614;
  wire  _T_1025 = _T_114 ? 1'h0 : _T_116;
  wire  _T_1026 = _T_112 ? 1'h0 : _T_1025;
  wire  _T_1027 = _T_110 ? 1'h0 : _T_1026;
  wire  _T_1028 = _T_108 ? 1'h0 : _T_1027;
  wire  _T_1029 = _T_106 ? 1'h0 : _T_1028;
  wire  _T_1030 = _T_104 ? 1'h0 : _T_1029;
  wire  _T_1031 = _T_102 ? 1'h0 : _T_1030;
  wire  _T_1032 = _T_100 ? 1'h0 : _T_1031;
  wire  _T_1033 = _T_98 ? 1'h0 : _T_1032;
  wire  _T_1034 = _T_96 ? 1'h0 : _T_1033;
  wire  _T_1035 = _T_94 ? 1'h0 : _T_1034;
  wire  _T_1036 = _T_92 ? 1'h0 : _T_1035;
  wire  _T_1037 = _T_90 ? 1'h0 : _T_1036;
  wire  _T_1038 = _T_88 ? 1'h0 : _T_1037;
  wire  _T_1039 = _T_86 ? 1'h0 : _T_1038;
  wire  _T_1040 = _T_84 ? 1'h0 : _T_1039;
  wire  _T_1041 = _T_82 ? 1'h0 : _T_1040;
  wire  _T_1042 = _T_80 ? 1'h0 : _T_1041;
  wire  _T_1043 = _T_78 ? 1'h0 : _T_1042;
  wire  _T_1044 = _T_76 ? 1'h0 : _T_1043;
  wire  _T_1045 = _T_74 ? 1'h0 : _T_1044;
  wire  _T_1046 = _T_72 ? 1'h0 : _T_1045;
  wire  _T_1047 = _T_70 ? 1'h0 : _T_1046;
  wire  _T_1048 = _T_68 ? 1'h0 : _T_1047;
  wire  _T_1049 = _T_66 ? 1'h0 : _T_1048;
  wire  _T_1050 = _T_64 ? 1'h0 : _T_1049;
  wire  _T_1051 = _T_62 ? 1'h0 : _T_1050;
  wire  _T_1052 = _T_60 ? 1'h0 : _T_1051;
  wire  _T_1053 = _T_58 ? 1'h0 : _T_1052;
  wire  _T_1054 = _T_56 ? 1'h0 : _T_1053;
  wire  _T_1055 = _T_54 ? 1'h0 : _T_1054;
  wire  _T_1056 = _T_52 ? 1'h0 : _T_1055;
  wire  _T_1057 = _T_50 ? 1'h0 : _T_1056;
  wire  _T_1058 = _T_48 ? 1'h0 : _T_1057;
  wire  _T_1059 = _T_46 ? 1'h0 : _T_1058;
  wire  _T_1060 = _T_44 ? 1'h0 : _T_1059;
  wire  _T_1061 = _T_42 ? 1'h0 : _T_1060;
  wire  _T_1062 = _T_40 ? 1'h0 : _T_1061;
  wire  c0_8 = _T_38 ? 1'h0 : _T_1062;
  wire  _T_1088 = _T_116 ? 1'h0 : _T_118;
  wire  _T_1089 = _T_114 ? 1'h0 : _T_1088;
  wire  _T_1090 = _T_112 ? 1'h0 : _T_1089;
  wire  _T_1091 = _T_110 ? 1'h0 : _T_1090;
  wire  _T_1092 = _T_108 ? 1'h0 : _T_1091;
  wire  _T_1093 = _T_106 ? 1'h0 : _T_1092;
  wire  _T_1094 = _T_104 ? 1'h0 : _T_1093;
  wire  _T_1095 = _T_102 ? 1'h0 : _T_1094;
  wire  _T_1096 = _T_100 ? 1'h0 : _T_1095;
  wire  _T_1097 = _T_98 ? 1'h0 : _T_1096;
  wire  _T_1098 = _T_96 ? 1'h0 : _T_1097;
  wire  _T_1099 = _T_94 ? 1'h0 : _T_1098;
  wire  _T_1100 = _T_92 ? 1'h0 : _T_1099;
  wire  _T_1101 = _T_90 ? 1'h0 : _T_1100;
  wire  _T_1102 = _T_88 ? 1'h0 : _T_1101;
  wire  _T_1103 = _T_86 ? 1'h0 : _T_1102;
  wire  _T_1104 = _T_84 ? 1'h0 : _T_1103;
  wire  _T_1105 = _T_82 ? 1'h0 : _T_1104;
  wire  _T_1106 = _T_80 ? 1'h0 : _T_1105;
  wire  _T_1107 = _T_78 ? 1'h0 : _T_1106;
  wire  _T_1108 = _T_76 ? 1'h0 : _T_1107;
  wire  _T_1109 = _T_74 ? 1'h0 : _T_1108;
  wire  _T_1110 = _T_72 ? 1'h0 : _T_1109;
  wire  _T_1111 = _T_70 ? 1'h0 : _T_1110;
  wire  _T_1112 = _T_68 ? 1'h0 : _T_1111;
  wire  _T_1113 = _T_66 ? 1'h0 : _T_1112;
  wire  _T_1114 = _T_64 ? 1'h0 : _T_1113;
  wire  _T_1115 = _T_62 ? 1'h0 : _T_1114;
  wire  _T_1116 = _T_60 ? 1'h0 : _T_1115;
  wire  _T_1117 = _T_58 ? 1'h0 : _T_1116;
  wire  _T_1118 = _T_56 ? 1'h0 : _T_1117;
  wire  _T_1119 = _T_54 ? 1'h0 : _T_1118;
  wire  _T_1120 = _T_52 ? 1'h0 : _T_1119;
  wire  _T_1121 = _T_50 ? 1'h0 : _T_1120;
  wire  _T_1122 = _T_48 ? 1'h0 : _T_1121;
  wire  _T_1123 = _T_46 ? 1'h0 : _T_1122;
  wire  _T_1124 = _T_44 ? 1'h0 : _T_1123;
  wire  _T_1125 = _T_42 ? 1'h0 : _T_1124;
  wire  _T_1126 = _T_40 ? 1'h0 : _T_1125;
  wire  c0_9 = _T_38 ? 1'h0 : _T_1126;
  wire [28:0] pa_lo_4 = EXVA[28:0];
  wire [31:0] _pa_T_6 = {csrs_27_PSEG,pa_lo_4};
  wire [31:0] _pa_T_7 = {csrs_28_PSEG,pa_lo_4};
  wire [19:0] _foundTLB_T_1197 = tlbHit_0_1 ? tlb_0_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1198 = tlbHit_1_1 ? tlb_1_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1199 = tlbHit_2_1 ? tlb_2_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1200 = tlbHit_3_1 ? tlb_3_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1201 = tlbHit_4_1 ? tlb_4_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1202 = tlbHit_5_1 ? tlb_5_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1203 = tlbHit_6_1 ? tlb_6_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1204 = tlbHit_7_1 ? tlb_7_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1205 = tlbHit_8_1 ? tlb_8_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1206 = tlbHit_9_1 ? tlb_9_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1207 = tlbHit_10_1 ? tlb_10_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1208 = tlbHit_11_1 ? tlb_11_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1209 = tlbHit_12_1 ? tlb_12_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1210 = tlbHit_13_1 ? tlb_13_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1211 = tlbHit_14_1 ? tlb_14_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1212 = tlbHit_15_1 ? tlb_15_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1213 = tlbHit_16_1 ? tlb_16_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1214 = tlbHit_17_1 ? tlb_17_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1215 = tlbHit_18_1 ? tlb_18_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1216 = tlbHit_19_1 ? tlb_19_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1217 = tlbHit_20_1 ? tlb_20_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1218 = tlbHit_21_1 ? tlb_21_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1219 = tlbHit_22_1 ? tlb_22_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1220 = tlbHit_23_1 ? tlb_23_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1221 = tlbHit_24_1 ? tlb_24_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1222 = tlbHit_25_1 ? tlb_25_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1223 = tlbHit_26_1 ? tlb_26_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1224 = tlbHit_27_1 ? tlb_27_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1225 = tlbHit_28_1 ? tlb_28_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1226 = tlbHit_29_1 ? tlb_29_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1227 = tlbHit_30_1 ? tlb_30_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1228 = tlbHit_31_1 ? tlb_31_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1229 = _foundTLB_T_1197 | _foundTLB_T_1198;
  wire [19:0] _foundTLB_T_1230 = _foundTLB_T_1229 | _foundTLB_T_1199;
  wire [19:0] _foundTLB_T_1231 = _foundTLB_T_1230 | _foundTLB_T_1200;
  wire [19:0] _foundTLB_T_1232 = _foundTLB_T_1231 | _foundTLB_T_1201;
  wire [19:0] _foundTLB_T_1233 = _foundTLB_T_1232 | _foundTLB_T_1202;
  wire [19:0] _foundTLB_T_1234 = _foundTLB_T_1233 | _foundTLB_T_1203;
  wire [19:0] _foundTLB_T_1235 = _foundTLB_T_1234 | _foundTLB_T_1204;
  wire [19:0] _foundTLB_T_1236 = _foundTLB_T_1235 | _foundTLB_T_1205;
  wire [19:0] _foundTLB_T_1237 = _foundTLB_T_1236 | _foundTLB_T_1206;
  wire [19:0] _foundTLB_T_1238 = _foundTLB_T_1237 | _foundTLB_T_1207;
  wire [19:0] _foundTLB_T_1239 = _foundTLB_T_1238 | _foundTLB_T_1208;
  wire [19:0] _foundTLB_T_1240 = _foundTLB_T_1239 | _foundTLB_T_1209;
  wire [19:0] _foundTLB_T_1241 = _foundTLB_T_1240 | _foundTLB_T_1210;
  wire [19:0] _foundTLB_T_1242 = _foundTLB_T_1241 | _foundTLB_T_1211;
  wire [19:0] _foundTLB_T_1243 = _foundTLB_T_1242 | _foundTLB_T_1212;
  wire [19:0] _foundTLB_T_1244 = _foundTLB_T_1243 | _foundTLB_T_1213;
  wire [19:0] _foundTLB_T_1245 = _foundTLB_T_1244 | _foundTLB_T_1214;
  wire [19:0] _foundTLB_T_1246 = _foundTLB_T_1245 | _foundTLB_T_1215;
  wire [19:0] _foundTLB_T_1247 = _foundTLB_T_1246 | _foundTLB_T_1216;
  wire [19:0] _foundTLB_T_1248 = _foundTLB_T_1247 | _foundTLB_T_1217;
  wire [19:0] _foundTLB_T_1249 = _foundTLB_T_1248 | _foundTLB_T_1218;
  wire [19:0] _foundTLB_T_1250 = _foundTLB_T_1249 | _foundTLB_T_1219;
  wire [19:0] _foundTLB_T_1251 = _foundTLB_T_1250 | _foundTLB_T_1220;
  wire [19:0] _foundTLB_T_1252 = _foundTLB_T_1251 | _foundTLB_T_1221;
  wire [19:0] _foundTLB_T_1253 = _foundTLB_T_1252 | _foundTLB_T_1222;
  wire [19:0] _foundTLB_T_1254 = _foundTLB_T_1253 | _foundTLB_T_1223;
  wire [19:0] _foundTLB_T_1255 = _foundTLB_T_1254 | _foundTLB_T_1224;
  wire [19:0] _foundTLB_T_1256 = _foundTLB_T_1255 | _foundTLB_T_1225;
  wire [19:0] _foundTLB_T_1257 = _foundTLB_T_1256 | _foundTLB_T_1226;
  wire [19:0] _foundTLB_T_1258 = _foundTLB_T_1257 | _foundTLB_T_1227;
  wire [19:0] foundTLB_1_P1_PPN = _foundTLB_T_1258 | _foundTLB_T_1228;
  wire [19:0] _foundTLB_T_1512 = tlbHit_0_1 ? tlb_0_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1513 = tlbHit_1_1 ? tlb_1_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1514 = tlbHit_2_1 ? tlb_2_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1515 = tlbHit_3_1 ? tlb_3_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1516 = tlbHit_4_1 ? tlb_4_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1517 = tlbHit_5_1 ? tlb_5_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1518 = tlbHit_6_1 ? tlb_6_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1519 = tlbHit_7_1 ? tlb_7_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1520 = tlbHit_8_1 ? tlb_8_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1521 = tlbHit_9_1 ? tlb_9_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1522 = tlbHit_10_1 ? tlb_10_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1523 = tlbHit_11_1 ? tlb_11_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1524 = tlbHit_12_1 ? tlb_12_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1525 = tlbHit_13_1 ? tlb_13_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1526 = tlbHit_14_1 ? tlb_14_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1527 = tlbHit_15_1 ? tlb_15_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1528 = tlbHit_16_1 ? tlb_16_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1529 = tlbHit_17_1 ? tlb_17_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1530 = tlbHit_18_1 ? tlb_18_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1531 = tlbHit_19_1 ? tlb_19_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1532 = tlbHit_20_1 ? tlb_20_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1533 = tlbHit_21_1 ? tlb_21_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1534 = tlbHit_22_1 ? tlb_22_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1535 = tlbHit_23_1 ? tlb_23_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1536 = tlbHit_24_1 ? tlb_24_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1537 = tlbHit_25_1 ? tlb_25_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1538 = tlbHit_26_1 ? tlb_26_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1539 = tlbHit_27_1 ? tlb_27_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1540 = tlbHit_28_1 ? tlb_28_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1541 = tlbHit_29_1 ? tlb_29_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1542 = tlbHit_30_1 ? tlb_30_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1543 = tlbHit_31_1 ? tlb_31_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_1544 = _foundTLB_T_1512 | _foundTLB_T_1513;
  wire [19:0] _foundTLB_T_1545 = _foundTLB_T_1544 | _foundTLB_T_1514;
  wire [19:0] _foundTLB_T_1546 = _foundTLB_T_1545 | _foundTLB_T_1515;
  wire [19:0] _foundTLB_T_1547 = _foundTLB_T_1546 | _foundTLB_T_1516;
  wire [19:0] _foundTLB_T_1548 = _foundTLB_T_1547 | _foundTLB_T_1517;
  wire [19:0] _foundTLB_T_1549 = _foundTLB_T_1548 | _foundTLB_T_1518;
  wire [19:0] _foundTLB_T_1550 = _foundTLB_T_1549 | _foundTLB_T_1519;
  wire [19:0] _foundTLB_T_1551 = _foundTLB_T_1550 | _foundTLB_T_1520;
  wire [19:0] _foundTLB_T_1552 = _foundTLB_T_1551 | _foundTLB_T_1521;
  wire [19:0] _foundTLB_T_1553 = _foundTLB_T_1552 | _foundTLB_T_1522;
  wire [19:0] _foundTLB_T_1554 = _foundTLB_T_1553 | _foundTLB_T_1523;
  wire [19:0] _foundTLB_T_1555 = _foundTLB_T_1554 | _foundTLB_T_1524;
  wire [19:0] _foundTLB_T_1556 = _foundTLB_T_1555 | _foundTLB_T_1525;
  wire [19:0] _foundTLB_T_1557 = _foundTLB_T_1556 | _foundTLB_T_1526;
  wire [19:0] _foundTLB_T_1558 = _foundTLB_T_1557 | _foundTLB_T_1527;
  wire [19:0] _foundTLB_T_1559 = _foundTLB_T_1558 | _foundTLB_T_1528;
  wire [19:0] _foundTLB_T_1560 = _foundTLB_T_1559 | _foundTLB_T_1529;
  wire [19:0] _foundTLB_T_1561 = _foundTLB_T_1560 | _foundTLB_T_1530;
  wire [19:0] _foundTLB_T_1562 = _foundTLB_T_1561 | _foundTLB_T_1531;
  wire [19:0] _foundTLB_T_1563 = _foundTLB_T_1562 | _foundTLB_T_1532;
  wire [19:0] _foundTLB_T_1564 = _foundTLB_T_1563 | _foundTLB_T_1533;
  wire [19:0] _foundTLB_T_1565 = _foundTLB_T_1564 | _foundTLB_T_1534;
  wire [19:0] _foundTLB_T_1566 = _foundTLB_T_1565 | _foundTLB_T_1535;
  wire [19:0] _foundTLB_T_1567 = _foundTLB_T_1566 | _foundTLB_T_1536;
  wire [19:0] _foundTLB_T_1568 = _foundTLB_T_1567 | _foundTLB_T_1537;
  wire [19:0] _foundTLB_T_1569 = _foundTLB_T_1568 | _foundTLB_T_1538;
  wire [19:0] _foundTLB_T_1570 = _foundTLB_T_1569 | _foundTLB_T_1539;
  wire [19:0] _foundTLB_T_1571 = _foundTLB_T_1570 | _foundTLB_T_1540;
  wire [19:0] _foundTLB_T_1572 = _foundTLB_T_1571 | _foundTLB_T_1541;
  wire [19:0] _foundTLB_T_1573 = _foundTLB_T_1572 | _foundTLB_T_1542;
  wire [19:0] foundTLB_1_P0_PPN = _foundTLB_T_1573 | _foundTLB_T_1543;
  wire [19:0] foundP_1_PPN = oddPG_1 ? foundTLB_1_P1_PPN : foundTLB_1_P0_PPN;
  wire [11:0] pa_lo_6 = EXVA[11:0];
  wire [31:0] _pa_T_9 = {foundP_1_PPN,pa_lo_6};
  wire [9:0] pa_hi_1 = foundP_1_PPN[19:10];
  wire [11:0] pa_lo_7 = EXVA[21:10];
  wire [21:0] _pa_T_10 = {pa_hi_1,pa_lo_7};
  wire [31:0] _pa_T_11 = _oddPG_T_3 ? _pa_T_9 : {{10'd0}, _pa_T_10};
  wire [31:0] _GEN_68 = EXVA[31:29] == csrs_28_VSEG & (csrs_28_PLV0 & _T_11 | csrs_28_PLV3 & _T_13) ? _pa_T_7 : _pa_T_11
    ;
  wire [31:0] pa_1 = EXVA[31:29] == csrs_27_VSEG & (csrs_27_PLV0 & crmd_PLV == 2'h0 | csrs_27_PLV3 & crmd_PLV == 2'h3)
     ? _pa_T_6 : _GEN_68;
  wire [3:0] _GEN_81 = 2'h1 == c0_3[2:1] ? 4'h3 : 4'h1;
  wire [3:0] _GEN_82 = 2'h2 == c0_3[2:1] ? 4'hf : _GEN_81;
  wire [3:0] _GEN_83 = 2'h3 == c0_3[2:1] ? 4'h0 : _GEN_82;
  wire [6:0] _GEN_4320 = {{3'd0}, _GEN_83};
  wire [6:0] memMask = _GEN_4320 << aluOut[1:0];
  wire  _GEN_88 = pme_1 & c0_2[0] ? c0_12 : 1'h1;
  wire  _GEN_92 = ppi_1 ? c0_12 : _GEN_88;
  wire  _GEN_98 = invalid_1 ? c0_12 : _GEN_92;
  wire  _GEN_105 = miss_1 ? c0_12 : _GEN_98;
  wire  _GEN_107 = crmd_DA | _GEN_105;
  wire  _GEN_115 = memADEM ? c0_12 : _GEN_107;
  wire  _GEN_124 = memALE ? c0_12 : _GEN_115;
  wire  _GEN_131 = c0_3 == 3'h7 | c0_11 & d[4:3] != 2'h2 | _GEN_124;
  wire  _GEN_145 = ID_OK & _GEN_131;
  wire  mem_OK = dStallReg | _GEN_145;
  wire  _GEN_89 = pme_1 & c0_2[0] & c0_12;
  wire  _GEN_93 = ppi_1 ? c0_12 : _GEN_89;
  wire  _GEN_99 = invalid_1 ? c0_12 : _GEN_93;
  wire  _GEN_106 = miss_1 ? c0_12 : _GEN_99;
  wire  _GEN_113 = crmd_DA ? c0_12 : _GEN_106;
  wire  _GEN_121 = memADEM ? c0_12 : _GEN_113;
  wire  _GEN_130 = memALE ? c0_12 : _GEN_121;
  wire  _GEN_139 = c0_3 == 3'h7 | c0_11 & d[4:3] != 2'h2 ? c0_12 : _GEN_130;
  wire  _GEN_153 = ID_OK ? _GEN_139 : c0_12;
  wire  preldNop = dStallReg ? c0_12 : _GEN_153;
  wire  _io_data_req_bits_wen_T_1 = c0_2 == 2'h3;
  wire [6:0] _io_data_req_bits_wen_T_4 = c0_2 == 2'h1 | c0_2 == 2'h3 & csrs_25_ROLLB ? memMask : 7'h0;
  wire [4:0] _io_data_req_bits_wdata_T_1 = {aluOut[1:0], 3'h0};
  wire [62:0] _GEN_4321 = {{31'd0}, rkd};
  wire [62:0] _io_data_req_bits_wdata_T_2 = _GEN_4321 << _io_data_req_bits_wdata_T_1;
  wire [31:0] shiftData = io_data_resp_bits >> _io_data_req_bits_wdata_T_1;
  wire  _extendData_T = c0_3 == 3'h0;
  wire [23:0] extendData_hi = shiftData[7] ? 24'hffffff : 24'h0;
  wire [7:0] extendData_lo = shiftData[7:0];
  wire [31:0] _extendData_T_3 = {extendData_hi,extendData_lo};
  wire  _extendData_T_4 = c0_3 == 3'h1;
  wire [31:0] _extendData_T_5 = {24'h0,extendData_lo};
  wire  _extendData_T_6 = c0_3 == 3'h2;
  wire [15:0] extendData_hi_1 = shiftData[15] ? 16'hffff : 16'h0;
  wire [15:0] extendData_lo_2 = shiftData[15:0];
  wire [31:0] _extendData_T_9 = {extendData_hi_1,extendData_lo_2};
  wire  _extendData_T_10 = c0_3 == 3'h3;
  wire [31:0] _extendData_T_11 = {16'h0,extendData_lo_2};
  wire  _extendData_T_12 = c0_3 == 3'h4;
  wire [31:0] _extendData_T_13 = _extendData_T ? _extendData_T_3 : 32'h0;
  wire [31:0] _extendData_T_14 = _extendData_T_4 ? _extendData_T_5 : 32'h0;
  wire [31:0] _extendData_T_15 = _extendData_T_6 ? _extendData_T_9 : 32'h0;
  wire [31:0] _extendData_T_16 = _extendData_T_10 ? _extendData_T_11 : 32'h0;
  wire [31:0] _extendData_T_17 = _extendData_T_12 ? shiftData : 32'h0;
  wire [31:0] _extendData_T_18 = _extendData_T_13 | _extendData_T_14;
  wire [31:0] _extendData_T_19 = _extendData_T_18 | _extendData_T_15;
  wire [31:0] _extendData_T_20 = _extendData_T_19 | _extendData_T_16;
  wire [31:0] extendData = _extendData_T_20 | _extendData_T_17;
  wire  _GEN_140 = c0_2 == 2'h2 & mem_OK | csrs_25_ROLLB;
  wire  _GEN_141 = _io_data_req_bits_wen_T_1 & mem_OK ? 1'h0 : _GEN_140;
  wire [18:0] _GEN_142 = ~ALE & ~ADEM ? aluOut[31:13] : _GEN_50;
  wire [31:0] _GEN_143 = ~mem_OK ? aluOut : _GEN_49;
  wire [18:0] _GEN_144 = ~mem_OK ? _GEN_142 : _GEN_50;
  wire  _GEN_154 = ID_OK ? _GEN_141 : csrs_25_ROLLB;
  wire [31:0] _GEN_155 = ID_OK ? _GEN_143 : _GEN_49;
  wire [18:0] _GEN_156 = ID_OK ? _GEN_144 : _GEN_50;
  wire  _GEN_166 = dStallReg ? csrs_25_ROLLB : _GEN_154;
  wire [31:0] _GEN_167 = dStallReg ? _GEN_49 : _GEN_155;
  wire [18:0] _GEN_168 = dStallReg ? _GEN_50 : _GEN_156;
  wire  dStall = ~io_data_resp_valid & (io_data_req_valid | dStallReg);
  wire  _csrRD_T = 14'h0 == SI14_lo;
  wire [8:0] _csrRD_T_1 = {crmd_DATM,crmd_DATF,crmd_PG,crmd_DA,crmd_IE,crmd_PLV};
  wire  _csrRD_T_2 = 14'h1 == SI14_lo;
  wire [2:0] _csrRD_T_3 = {csrs_1_PIE,csrs_1_PPLV};
  wire  _csrRD_T_4 = 14'h2 == SI14_lo;
  wire  _csrRD_T_5 = 14'h4 == SI14_lo;
  wire  _csrRD_T_6 = 14'h5 == SI14_lo;
  wire [7:0] csrRD_lo_1 = {csrs_4_IS_7,csrs_4_IS_6,csrs_4_IS_5,csrs_4_IS_4,csrs_4_IS_3,csrs_4_IS_2,csrs_4_IS_1,
    csrs_4_IS_0};
  wire [30:0] _csrRD_T_7 = {csrs_4_EsubCode,csrs_4_Ecode,3'h0,csrs_4_IS_12,csrs_4_IS_11,1'h0,csrs_4_IS_9,csrs_4_IS_8,
    csrRD_lo_1};
  wire  _csrRD_T_8 = 14'h6 == SI14_lo;
  wire  _csrRD_T_9 = 14'h7 == SI14_lo;
  wire  _csrRD_T_10 = 14'hc == SI14_lo;
  wire [31:0] _csrRD_T_11 = {csrs_7_VA,6'h0};
  wire  _csrRD_T_12 = 14'h10 == SI14_lo;
  wire [31:0] _csrRD_T_13 = {csrs_8_NE,1'h0,csrs_8_PS,19'h0,csrs_8_Index};
  wire  _csrRD_T_14 = 14'h11 == SI14_lo;
  wire  _csrRD_T_16 = 14'h12 == SI14_lo;
  wire [31:0] _csrRD_T_17 = {csrs_10_PPN,1'h0,csrs_10_G,csrs_10_MAT,csrs_10_PLV,csrs_10_D,csrs_10_V};
  wire  _csrRD_T_18 = 14'h13 == SI14_lo;
  wire [31:0] _csrRD_T_19 = {csrs_11_PPN,1'h0,csrs_11_G,csrs_11_MAT,csrs_11_PLV,csrs_11_D,csrs_11_V};
  wire  _csrRD_T_20 = 14'h18 == SI14_lo;
  wire [23:0] _csrRD_T_21 = {14'h280,asid_ASID};
  wire  _csrRD_T_22 = 14'h19 == SI14_lo;
  wire [31:0] _csrRD_T_23 = {csrs_13_Base,12'h0};
  wire  _csrRD_T_24 = 14'h1a == SI14_lo;
  wire [31:0] _csrRD_T_25 = {csrs_14_Base,12'h0};
  wire  _csrRD_T_26 = 14'h1b == SI14_lo;
  wire [31:0] _csrRD_T_30 = badv_VAddr[31] ? _csrRD_T_25 : _csrRD_T_23;
  wire  _csrRD_T_32 = 14'h30 == SI14_lo;
  wire  _csrRD_T_33 = 14'h31 == SI14_lo;
  wire  _csrRD_T_34 = 14'h32 == SI14_lo;
  wire  _csrRD_T_35 = 14'h33 == SI14_lo;
  wire  _csrRD_T_36 = 14'h40 == SI14_lo;
  wire  _csrRD_T_37 = 14'h41 == SI14_lo;
  wire [31:0] _csrRD_T_38 = {csrs_22_InitVal,csrs_22_Periodic,csrs_22_En};
  wire  _csrRD_T_39 = 14'h42 == SI14_lo;
  wire  _csrRD_T_40 = 14'h44 == SI14_lo;
  wire  _csrRD_T_41 = 14'h60 == SI14_lo;
  wire [2:0] _csrRD_T_42 = {csrs_25_KLO,1'h0,csrs_25_ROLLB};
  wire  _csrRD_T_43 = 14'h88 == SI14_lo;
  wire [31:0] _csrRD_T_44 = {csrs_26_PA,6'h0};
  wire  _csrRD_T_45 = 14'h180 == SI14_lo;
  wire [31:0] _csrRD_T_46 = {csrs_27_VSEG,1'h0,csrs_27_PSEG,19'h0,csrs_27_MAT,csrs_27_PLV3,2'h0,csrs_27_PLV0};
  wire  _csrRD_T_47 = 14'h181 == SI14_lo;
  wire [31:0] _csrRD_T_48 = {csrs_28_VSEG,1'h0,csrs_28_PSEG,19'h0,csrs_28_MAT,csrs_28_PLV3,2'h0,csrs_28_PLV0};
  wire [8:0] _csrRD_T_49 = _csrRD_T ? _csrRD_T_1 : 9'h0;
  wire [2:0] _csrRD_T_50 = _csrRD_T_2 ? _csrRD_T_3 : 3'h0;
  wire  _csrRD_T_51 = _csrRD_T_4 & csrs_2_FPE;
  wire [12:0] _csrRD_T_52 = _csrRD_T_5 ? csrs_3_LIE : 13'h0;
  wire [30:0] _csrRD_T_53 = _csrRD_T_6 ? _csrRD_T_7 : 31'h0;
  wire [31:0] _csrRD_T_54 = _csrRD_T_8 ? csrs_5_PC : 32'h0;
  wire [31:0] _csrRD_T_55 = _csrRD_T_9 ? badv_VAddr : 32'h0;
  wire [31:0] _csrRD_T_56 = _csrRD_T_10 ? _csrRD_T_11 : 32'h0;
  wire [31:0] _csrRD_T_57 = _csrRD_T_12 ? _csrRD_T_13 : 32'h0;
  wire [31:0] _csrRD_T_58 = _csrRD_T_14 ? _EXVA_T_2 : 32'h0;
  wire [31:0] _csrRD_T_59 = _csrRD_T_16 ? _csrRD_T_17 : 32'h0;
  wire [31:0] _csrRD_T_60 = _csrRD_T_18 ? _csrRD_T_19 : 32'h0;
  wire [23:0] _csrRD_T_61 = _csrRD_T_20 ? _csrRD_T_21 : 24'h0;
  wire [31:0] _csrRD_T_62 = _csrRD_T_22 ? _csrRD_T_23 : 32'h0;
  wire [31:0] _csrRD_T_63 = _csrRD_T_24 ? _csrRD_T_25 : 32'h0;
  wire [31:0] _csrRD_T_64 = _csrRD_T_26 ? _csrRD_T_30 : 32'h0;
  wire [31:0] _csrRD_T_66 = _csrRD_T_32 ? csrs_17_Data : 32'h0;
  wire [31:0] _csrRD_T_67 = _csrRD_T_33 ? csrs_18_Data : 32'h0;
  wire [31:0] _csrRD_T_68 = _csrRD_T_34 ? csrs_19_Data : 32'h0;
  wire [31:0] _csrRD_T_69 = _csrRD_T_35 ? csrs_20_Data : 32'h0;
  wire [31:0] _csrRD_T_70 = _csrRD_T_36 ? csrs_21_TID : 32'h0;
  wire [31:0] _csrRD_T_71 = _csrRD_T_37 ? _csrRD_T_38 : 32'h0;
  wire [31:0] _csrRD_T_72 = _csrRD_T_39 ? csrs_23_TimeVal : 32'h0;
  wire [2:0] _csrRD_T_74 = _csrRD_T_41 ? _csrRD_T_42 : 3'h0;
  wire [31:0] _csrRD_T_75 = _csrRD_T_43 ? _csrRD_T_44 : 32'h0;
  wire [31:0] _csrRD_T_76 = _csrRD_T_45 ? _csrRD_T_46 : 32'h0;
  wire [31:0] _csrRD_T_77 = _csrRD_T_47 ? _csrRD_T_48 : 32'h0;
  wire [8:0] _GEN_4322 = {{6'd0}, _csrRD_T_50};
  wire [8:0] _csrRD_T_78 = _csrRD_T_49 | _GEN_4322;
  wire [8:0] _GEN_4323 = {{8'd0}, _csrRD_T_51};
  wire [8:0] _csrRD_T_79 = _csrRD_T_78 | _GEN_4323;
  wire [12:0] _GEN_4324 = {{4'd0}, _csrRD_T_79};
  wire [12:0] _csrRD_T_80 = _GEN_4324 | _csrRD_T_52;
  wire [30:0] _GEN_4325 = {{18'd0}, _csrRD_T_80};
  wire [30:0] _csrRD_T_81 = _GEN_4325 | _csrRD_T_53;
  wire [31:0] _GEN_4326 = {{1'd0}, _csrRD_T_81};
  wire [31:0] _csrRD_T_82 = _GEN_4326 | _csrRD_T_54;
  wire [31:0] _csrRD_T_83 = _csrRD_T_82 | _csrRD_T_55;
  wire [31:0] _csrRD_T_84 = _csrRD_T_83 | _csrRD_T_56;
  wire [31:0] _csrRD_T_85 = _csrRD_T_84 | _csrRD_T_57;
  wire [31:0] _csrRD_T_86 = _csrRD_T_85 | _csrRD_T_58;
  wire [31:0] _csrRD_T_87 = _csrRD_T_86 | _csrRD_T_59;
  wire [31:0] _csrRD_T_88 = _csrRD_T_87 | _csrRD_T_60;
  wire [31:0] _GEN_4327 = {{8'd0}, _csrRD_T_61};
  wire [31:0] _csrRD_T_89 = _csrRD_T_88 | _GEN_4327;
  wire [31:0] _csrRD_T_90 = _csrRD_T_89 | _csrRD_T_62;
  wire [31:0] _csrRD_T_91 = _csrRD_T_90 | _csrRD_T_63;
  wire [31:0] _csrRD_T_92 = _csrRD_T_91 | _csrRD_T_64;
  wire [31:0] _csrRD_T_94 = _csrRD_T_92 | _csrRD_T_66;
  wire [31:0] _csrRD_T_95 = _csrRD_T_94 | _csrRD_T_67;
  wire [31:0] _csrRD_T_96 = _csrRD_T_95 | _csrRD_T_68;
  wire [31:0] _csrRD_T_97 = _csrRD_T_96 | _csrRD_T_69;
  wire [31:0] _csrRD_T_98 = _csrRD_T_97 | _csrRD_T_70;
  wire [31:0] _csrRD_T_99 = _csrRD_T_98 | _csrRD_T_71;
  wire [31:0] _csrRD_T_100 = _csrRD_T_99 | _csrRD_T_72;
  wire [31:0] _GEN_4328 = {{29'd0}, _csrRD_T_74};
  wire [31:0] _csrRD_T_102 = _csrRD_T_100 | _GEN_4328;
  wire [31:0] _csrRD_T_103 = _csrRD_T_102 | _csrRD_T_75;
  wire [31:0] _csrRD_T_104 = _csrRD_T_103 | _csrRD_T_76;
  wire [31:0] csrRD = _csrRD_T_104 | _csrRD_T_77;
  wire [31:0] csrMask = j == 5'h1 ? 32'hffffffff : rj;
  wire [31:0] _crmd_T = rkd & csrMask;
  wire [31:0] _crmd_T_2 = ~csrMask;
  wire [31:0] _GEN_4329 = {{23'd0}, _csrRD_T_1};
  wire [31:0] _crmd_T_3 = _GEN_4329 & _crmd_T_2;
  wire [31:0] _crmd_T_4 = _crmd_T | _crmd_T_3;
  wire [1:0] _GEN_169 = _csrRD_T ? _crmd_T_4[1:0] : crmd_PLV;
  wire  _GEN_170 = _csrRD_T ? _crmd_T_4[2] : crmd_IE;
  wire  _GEN_171 = _csrRD_T ? _crmd_T_4[3] : crmd_DA;
  wire  _GEN_172 = _csrRD_T ? _crmd_T_4[4] : crmd_PG;
  wire [31:0] _GEN_4330 = {{29'd0}, _csrRD_T_3};
  wire [31:0] _prmd_T_3 = _GEN_4330 & _crmd_T_2;
  wire [31:0] _prmd_T_4 = _crmd_T | _prmd_T_3;
  wire [1:0] _GEN_175 = _csrRD_T_2 ? _prmd_T_4[1:0] : csrs_1_PPLV;
  wire  _GEN_176 = _csrRD_T_2 ? _prmd_T_4[2] : csrs_1_PIE;
  wire [31:0] _GEN_4331 = {{31'd0}, csrs_2_FPE};
  wire [31:0] _euen_T_2 = _GEN_4331 & _crmd_T_2;
  wire [31:0] _euen_T_3 = _crmd_T | _euen_T_2;
  wire [31:0] _GEN_4332 = {{19'd0}, csrs_3_LIE};
  wire [31:0] _ectl_T_2 = _GEN_4332 & _crmd_T_2;
  wire [31:0] _ectl_T_3 = _crmd_T | _ectl_T_2;
  wire [31:0] _era_T_2 = csrs_5_PC & _crmd_T_2;
  wire [31:0] _era_T_3 = _crmd_T | _era_T_2;
  wire [31:0] _GEN_183 = _csrRD_T_8 ? _era_T_3 : csrs_5_PC;
  wire [31:0] _badv_T_2 = badv_VAddr & _crmd_T_2;
  wire [31:0] _badv_T_3 = _crmd_T | _badv_T_2;
  wire [25:0] _eentry_VA_T = rkd[31:6] & csrMask[31:6];
  wire [25:0] _eentry_VA_T_1 = ~csrMask[31:6];
  wire [25:0] _eentry_VA_T_2 = csrs_7_VA & _eentry_VA_T_1;
  wire [25:0] _eentry_VA_T_3 = _eentry_VA_T | _eentry_VA_T_2;
  wire [5:0] _tlbidx_PS_T = rkd[29:24] & csrMask[29:24];
  wire [5:0] _tlbidx_PS_T_1 = ~csrMask[29:24];
  wire [5:0] _tlbidx_PS_T_2 = csrs_8_PS & _tlbidx_PS_T_1;
  wire [5:0] _tlbidx_PS_T_3 = _tlbidx_PS_T | _tlbidx_PS_T_2;
  wire [4:0] _tlbidx_Index_T = rkd[4:0] & csrMask[4:0];
  wire [4:0] _tlbidx_Index_T_1 = ~csrMask[4:0];
  wire [4:0] _tlbidx_Index_T_2 = csrs_8_Index & _tlbidx_Index_T_1;
  wire [4:0] _tlbidx_Index_T_3 = _tlbidx_Index_T | _tlbidx_Index_T_2;
  wire  _GEN_186 = _csrRD_T_12 ? rkd[31] & csrMask[31] | csrs_8_NE & ~csrMask[31] : csrs_8_NE;
  wire [5:0] _GEN_187 = _csrRD_T_12 ? _tlbidx_PS_T_3 : csrs_8_PS;
  wire [4:0] _GEN_188 = _csrRD_T_12 ? _tlbidx_Index_T_3 : csrs_8_Index;
  wire [18:0] _tlbehi_VPPN_T_2 = rkd[31:13] & csrMask[31:13];
  wire [18:0] _tlbehi_VPPN_T_3 = ~csrMask[31:13];
  wire [18:0] _tlbehi_VPPN_T_4 = csrs_9_VPPN & _tlbehi_VPPN_T_3;
  wire [18:0] _tlbehi_VPPN_T_5 = _tlbehi_VPPN_T_2 | _tlbehi_VPPN_T_4;
  wire [18:0] _GEN_189 = _csrRD_T_14 ? _tlbehi_VPPN_T_5 : _GEN_168;
  wire [31:0] _tlbelo0_T_3 = _csrRD_T_17 & _crmd_T_2;
  wire [31:0] _tlbelo0_T_4 = _crmd_T | _tlbelo0_T_3;
  wire [23:0] _tlbelo0_PPN_T = rkd[31:8] & csrMask[31:8];
  wire [23:0] _tlbelo0_PPN_T_1 = ~csrMask[31:8];
  wire [23:0] _tlbelo0_PPN_T_2 = csrs_10_PPN & _tlbelo0_PPN_T_1;
  wire [23:0] _tlbelo0_PPN_T_3 = _tlbelo0_PPN_T | _tlbelo0_PPN_T_2;
  wire  _GEN_190 = _csrRD_T_16 ? _tlbelo0_T_4[0] : csrs_10_V;
  wire  _GEN_191 = _csrRD_T_16 ? _tlbelo0_T_4[1] : csrs_10_D;
  wire [1:0] _GEN_192 = _csrRD_T_16 ? _tlbelo0_T_4[3:2] : csrs_10_PLV;
  wire [1:0] _GEN_193 = _csrRD_T_16 ? _tlbelo0_T_4[5:4] : csrs_10_MAT;
  wire  _GEN_194 = _csrRD_T_16 ? _tlbelo0_T_4[6] : csrs_10_G;
  wire [23:0] _GEN_195 = _csrRD_T_16 ? _tlbelo0_PPN_T_3 : csrs_10_PPN;
  wire [31:0] _tlbelo1_T_3 = _csrRD_T_19 & _crmd_T_2;
  wire [31:0] _tlbelo1_T_4 = _crmd_T | _tlbelo1_T_3;
  wire [23:0] _tlbelo1_PPN_T_2 = csrs_11_PPN & _tlbelo0_PPN_T_1;
  wire [23:0] _tlbelo1_PPN_T_3 = _tlbelo0_PPN_T | _tlbelo1_PPN_T_2;
  wire  _GEN_196 = _csrRD_T_18 ? _tlbelo1_T_4[0] : csrs_11_V;
  wire  _GEN_197 = _csrRD_T_18 ? _tlbelo1_T_4[1] : csrs_11_D;
  wire [1:0] _GEN_198 = _csrRD_T_18 ? _tlbelo1_T_4[3:2] : csrs_11_PLV;
  wire [1:0] _GEN_199 = _csrRD_T_18 ? _tlbelo1_T_4[5:4] : csrs_11_MAT;
  wire  _GEN_200 = _csrRD_T_18 ? _tlbelo1_T_4[6] : csrs_11_G;
  wire [23:0] _GEN_201 = _csrRD_T_18 ? _tlbelo1_PPN_T_3 : csrs_11_PPN;
  wire [9:0] _asid_ASID_T = rkd[9:0] & csrMask[9:0];
  wire [9:0] _asid_ASID_T_1 = ~csrMask[9:0];
  wire [9:0] _asid_ASID_T_2 = asid_ASID & _asid_ASID_T_1;
  wire [9:0] _asid_ASID_T_3 = _asid_ASID_T | _asid_ASID_T_2;
  wire [9:0] _GEN_202 = _csrRD_T_20 ? _asid_ASID_T_3 : asid_ASID;
  wire [19:0] _pgdl_Base_T = rkd[31:12] & csrMask[31:12];
  wire [19:0] _pgdl_Base_T_1 = ~csrMask[31:12];
  wire [19:0] _pgdl_Base_T_2 = csrs_13_Base & _pgdl_Base_T_1;
  wire [19:0] _pgdl_Base_T_3 = _pgdl_Base_T | _pgdl_Base_T_2;
  wire [19:0] _pgdh_Base_T_2 = csrs_14_Base & _pgdl_Base_T_1;
  wire [19:0] _pgdh_Base_T_3 = _pgdl_Base_T | _pgdh_Base_T_2;
  wire [31:0] _save0_T_2 = csrs_17_Data & _crmd_T_2;
  wire [31:0] _save0_T_3 = _crmd_T | _save0_T_2;
  wire [31:0] _save1_T_2 = csrs_18_Data & _crmd_T_2;
  wire [31:0] _save1_T_3 = _crmd_T | _save1_T_2;
  wire [31:0] _save2_T_2 = csrs_19_Data & _crmd_T_2;
  wire [31:0] _save2_T_3 = _crmd_T | _save2_T_2;
  wire [31:0] _save3_T_2 = csrs_20_Data & _crmd_T_2;
  wire [31:0] _save3_T_3 = _crmd_T | _save3_T_2;
  wire [31:0] _tid_T_2 = csrs_21_TID & _crmd_T_2;
  wire [31:0] _tid_T_3 = _crmd_T | _tid_T_2;
  wire [31:0] _tcfg_T_3 = _csrRD_T_38 & _crmd_T_2;
  wire [31:0] _tcfg_T_4 = _crmd_T | _tcfg_T_3;
  wire [31:0] _T_1407 = rkd & 32'hfffffffc;
  wire [31:0] _tval_TimeVal_T_3 = _T_1407 & csrMask;
  wire [31:0] _tval_TimeVal_T_5 = csrs_23_TimeVal & _crmd_T_2;
  wire [31:0] _tval_TimeVal_T_6 = _tval_TimeVal_T_3 | _tval_TimeVal_T_5;
  wire  _T_1412 = rkd[0] & csrMask[0];
  wire  _GEN_216 = csrMask[2] ? rkd[2] : csrs_25_KLO;
  wire  _GEN_217 = csrMask[1] & rkd[1] ? 1'h0 : _GEN_166;
  wire  _GEN_219 = _csrRD_T_41 ? _GEN_217 : _GEN_166;
  wire [25:0] _tlbrentry_PA_T_2 = csrs_26_PA & _eentry_VA_T_1;
  wire [25:0] _tlbrentry_PA_T_3 = _eentry_VA_T | _tlbrentry_PA_T_2;
  wire [1:0] _dmw0_MAT_T = rkd[5:4] & csrMask[5:4];
  wire [1:0] _dmw0_MAT_T_1 = ~csrMask[5:4];
  wire [1:0] _dmw0_MAT_T_2 = csrs_27_MAT & _dmw0_MAT_T_1;
  wire [1:0] _dmw0_MAT_T_3 = _dmw0_MAT_T | _dmw0_MAT_T_2;
  wire [2:0] _dmw0_PSEG_T = rkd[27:25] & csrMask[27:25];
  wire [2:0] _dmw0_PSEG_T_1 = ~csrMask[27:25];
  wire [2:0] _dmw0_PSEG_T_2 = csrs_27_PSEG & _dmw0_PSEG_T_1;
  wire [2:0] _dmw0_PSEG_T_3 = _dmw0_PSEG_T | _dmw0_PSEG_T_2;
  wire [2:0] _dmw0_VSEG_T = rkd[31:29] & csrMask[31:29];
  wire [2:0] _dmw0_VSEG_T_1 = ~csrMask[31:29];
  wire [2:0] _dmw0_VSEG_T_2 = csrs_27_VSEG & _dmw0_VSEG_T_1;
  wire [2:0] _dmw0_VSEG_T_3 = _dmw0_VSEG_T | _dmw0_VSEG_T_2;
  wire [1:0] _dmw1_MAT_T_2 = csrs_28_MAT & _dmw0_MAT_T_1;
  wire [1:0] _dmw1_MAT_T_3 = _dmw0_MAT_T | _dmw1_MAT_T_2;
  wire [2:0] _dmw1_PSEG_T_2 = csrs_28_PSEG & _dmw0_PSEG_T_1;
  wire [2:0] _dmw1_PSEG_T_3 = _dmw0_PSEG_T | _dmw1_PSEG_T_2;
  wire [2:0] _dmw1_VSEG_T_2 = csrs_28_VSEG & _dmw0_VSEG_T_1;
  wire [2:0] _dmw1_VSEG_T_3 = _dmw0_VSEG_T | _dmw1_VSEG_T_2;
  wire [1:0] _GEN_231 = ID_OK & c0_4 & |csrMask ? _GEN_169 : crmd_PLV;
  wire  _GEN_232 = ID_OK & c0_4 & |csrMask ? _GEN_170 : crmd_IE;
  wire  _GEN_233 = ID_OK & c0_4 & |csrMask ? _GEN_171 : crmd_DA;
  wire  _GEN_234 = ID_OK & c0_4 & |csrMask ? _GEN_172 : crmd_PG;
  wire [1:0] _GEN_237 = ID_OK & c0_4 & |csrMask ? _GEN_175 : csrs_1_PPLV;
  wire  _GEN_238 = ID_OK & c0_4 & |csrMask ? _GEN_176 : csrs_1_PIE;
  wire [31:0] _GEN_243 = ID_OK & c0_4 & |csrMask ? _GEN_183 : csrs_5_PC;
  wire  _GEN_246 = ID_OK & c0_4 & |csrMask ? _GEN_186 : csrs_8_NE;
  wire [5:0] _GEN_247 = ID_OK & c0_4 & |csrMask ? _GEN_187 : csrs_8_PS;
  wire [4:0] _GEN_248 = ID_OK & c0_4 & |csrMask ? _GEN_188 : csrs_8_Index;
  wire [18:0] _GEN_249 = ID_OK & c0_4 & |csrMask ? _GEN_189 : _GEN_168;
  wire  _GEN_250 = ID_OK & c0_4 & |csrMask ? _GEN_190 : csrs_10_V;
  wire  _GEN_251 = ID_OK & c0_4 & |csrMask ? _GEN_191 : csrs_10_D;
  wire [1:0] _GEN_252 = ID_OK & c0_4 & |csrMask ? _GEN_192 : csrs_10_PLV;
  wire [1:0] _GEN_253 = ID_OK & c0_4 & |csrMask ? _GEN_193 : csrs_10_MAT;
  wire  _GEN_254 = ID_OK & c0_4 & |csrMask ? _GEN_194 : csrs_10_G;
  wire [23:0] _GEN_255 = ID_OK & c0_4 & |csrMask ? _GEN_195 : csrs_10_PPN;
  wire  _GEN_256 = ID_OK & c0_4 & |csrMask ? _GEN_196 : csrs_11_V;
  wire  _GEN_257 = ID_OK & c0_4 & |csrMask ? _GEN_197 : csrs_11_D;
  wire [1:0] _GEN_258 = ID_OK & c0_4 & |csrMask ? _GEN_198 : csrs_11_PLV;
  wire [1:0] _GEN_259 = ID_OK & c0_4 & |csrMask ? _GEN_199 : csrs_11_MAT;
  wire  _GEN_260 = ID_OK & c0_4 & |csrMask ? _GEN_200 : csrs_11_G;
  wire [23:0] _GEN_261 = ID_OK & c0_4 & |csrMask ? _GEN_201 : csrs_11_PPN;
  wire [9:0] _GEN_262 = ID_OK & c0_4 & |csrMask ? _GEN_202 : asid_ASID;
  wire  _GEN_276 = ID_OK & c0_4 & |csrMask ? _GEN_219 : _GEN_166;
  wire [4:0] _tlbidx_Index_T_5 = tlbHit_1_1 ? 5'h1 : 5'h0;
  wire [4:0] _tlbidx_Index_T_6 = tlbHit_2_1 ? 5'h2 : 5'h0;
  wire [4:0] _tlbidx_Index_T_7 = tlbHit_3_1 ? 5'h3 : 5'h0;
  wire [4:0] _tlbidx_Index_T_8 = tlbHit_4_1 ? 5'h4 : 5'h0;
  wire [4:0] _tlbidx_Index_T_9 = tlbHit_5_1 ? 5'h5 : 5'h0;
  wire [4:0] _tlbidx_Index_T_10 = tlbHit_6_1 ? 5'h6 : 5'h0;
  wire [4:0] _tlbidx_Index_T_11 = tlbHit_7_1 ? 5'h7 : 5'h0;
  wire [4:0] _tlbidx_Index_T_12 = tlbHit_8_1 ? 5'h8 : 5'h0;
  wire [4:0] _tlbidx_Index_T_13 = tlbHit_9_1 ? 5'h9 : 5'h0;
  wire [4:0] _tlbidx_Index_T_14 = tlbHit_10_1 ? 5'ha : 5'h0;
  wire [4:0] _tlbidx_Index_T_15 = tlbHit_11_1 ? 5'hb : 5'h0;
  wire [4:0] _tlbidx_Index_T_16 = tlbHit_12_1 ? 5'hc : 5'h0;
  wire [4:0] _tlbidx_Index_T_17 = tlbHit_13_1 ? 5'hd : 5'h0;
  wire [4:0] _tlbidx_Index_T_18 = tlbHit_14_1 ? 5'he : 5'h0;
  wire [4:0] _tlbidx_Index_T_19 = tlbHit_15_1 ? 5'hf : 5'h0;
  wire [4:0] _tlbidx_Index_T_20 = tlbHit_16_1 ? 5'h10 : 5'h0;
  wire [4:0] _tlbidx_Index_T_21 = tlbHit_17_1 ? 5'h11 : 5'h0;
  wire [4:0] _tlbidx_Index_T_22 = tlbHit_18_1 ? 5'h12 : 5'h0;
  wire [4:0] _tlbidx_Index_T_23 = tlbHit_19_1 ? 5'h13 : 5'h0;
  wire [4:0] _tlbidx_Index_T_24 = tlbHit_20_1 ? 5'h14 : 5'h0;
  wire [4:0] _tlbidx_Index_T_25 = tlbHit_21_1 ? 5'h15 : 5'h0;
  wire [4:0] _tlbidx_Index_T_26 = tlbHit_22_1 ? 5'h16 : 5'h0;
  wire [4:0] _tlbidx_Index_T_27 = tlbHit_23_1 ? 5'h17 : 5'h0;
  wire [4:0] _tlbidx_Index_T_28 = tlbHit_24_1 ? 5'h18 : 5'h0;
  wire [4:0] _tlbidx_Index_T_29 = tlbHit_25_1 ? 5'h19 : 5'h0;
  wire [4:0] _tlbidx_Index_T_30 = tlbHit_26_1 ? 5'h1a : 5'h0;
  wire [4:0] _tlbidx_Index_T_31 = tlbHit_27_1 ? 5'h1b : 5'h0;
  wire [4:0] _tlbidx_Index_T_32 = tlbHit_28_1 ? 5'h1c : 5'h0;
  wire [4:0] _tlbidx_Index_T_33 = tlbHit_29_1 ? 5'h1d : 5'h0;
  wire [4:0] _tlbidx_Index_T_34 = tlbHit_30_1 ? 5'h1e : 5'h0;
  wire [4:0] _tlbidx_Index_T_35 = tlbHit_31_1 ? 5'h1f : 5'h0;
  wire [4:0] _tlbidx_Index_T_37 = _tlbidx_Index_T_5 | _tlbidx_Index_T_6;
  wire [4:0] _tlbidx_Index_T_38 = _tlbidx_Index_T_37 | _tlbidx_Index_T_7;
  wire [4:0] _tlbidx_Index_T_39 = _tlbidx_Index_T_38 | _tlbidx_Index_T_8;
  wire [4:0] _tlbidx_Index_T_40 = _tlbidx_Index_T_39 | _tlbidx_Index_T_9;
  wire [4:0] _tlbidx_Index_T_41 = _tlbidx_Index_T_40 | _tlbidx_Index_T_10;
  wire [4:0] _tlbidx_Index_T_42 = _tlbidx_Index_T_41 | _tlbidx_Index_T_11;
  wire [4:0] _tlbidx_Index_T_43 = _tlbidx_Index_T_42 | _tlbidx_Index_T_12;
  wire [4:0] _tlbidx_Index_T_44 = _tlbidx_Index_T_43 | _tlbidx_Index_T_13;
  wire [4:0] _tlbidx_Index_T_45 = _tlbidx_Index_T_44 | _tlbidx_Index_T_14;
  wire [4:0] _tlbidx_Index_T_46 = _tlbidx_Index_T_45 | _tlbidx_Index_T_15;
  wire [4:0] _tlbidx_Index_T_47 = _tlbidx_Index_T_46 | _tlbidx_Index_T_16;
  wire [4:0] _tlbidx_Index_T_48 = _tlbidx_Index_T_47 | _tlbidx_Index_T_17;
  wire [4:0] _tlbidx_Index_T_49 = _tlbidx_Index_T_48 | _tlbidx_Index_T_18;
  wire [4:0] _tlbidx_Index_T_50 = _tlbidx_Index_T_49 | _tlbidx_Index_T_19;
  wire [4:0] _tlbidx_Index_T_51 = _tlbidx_Index_T_50 | _tlbidx_Index_T_20;
  wire [4:0] _tlbidx_Index_T_52 = _tlbidx_Index_T_51 | _tlbidx_Index_T_21;
  wire [4:0] _tlbidx_Index_T_53 = _tlbidx_Index_T_52 | _tlbidx_Index_T_22;
  wire [4:0] _tlbidx_Index_T_54 = _tlbidx_Index_T_53 | _tlbidx_Index_T_23;
  wire [4:0] _tlbidx_Index_T_55 = _tlbidx_Index_T_54 | _tlbidx_Index_T_24;
  wire [4:0] _tlbidx_Index_T_56 = _tlbidx_Index_T_55 | _tlbidx_Index_T_25;
  wire [4:0] _tlbidx_Index_T_57 = _tlbidx_Index_T_56 | _tlbidx_Index_T_26;
  wire [4:0] _tlbidx_Index_T_58 = _tlbidx_Index_T_57 | _tlbidx_Index_T_27;
  wire [4:0] _tlbidx_Index_T_59 = _tlbidx_Index_T_58 | _tlbidx_Index_T_28;
  wire [4:0] _tlbidx_Index_T_60 = _tlbidx_Index_T_59 | _tlbidx_Index_T_29;
  wire [4:0] _tlbidx_Index_T_61 = _tlbidx_Index_T_60 | _tlbidx_Index_T_30;
  wire [4:0] _tlbidx_Index_T_62 = _tlbidx_Index_T_61 | _tlbidx_Index_T_31;
  wire [4:0] _tlbidx_Index_T_63 = _tlbidx_Index_T_62 | _tlbidx_Index_T_32;
  wire [4:0] _tlbidx_Index_T_64 = _tlbidx_Index_T_63 | _tlbidx_Index_T_33;
  wire [4:0] _tlbidx_Index_T_65 = _tlbidx_Index_T_64 | _tlbidx_Index_T_34;
  wire [4:0] _tlbidx_Index_T_66 = _tlbidx_Index_T_65 | _tlbidx_Index_T_35;
  wire  _GEN_291 = 5'h1 == csrs_8_Index ? tlb_1_E : tlb_0_E;
  wire  _GEN_292 = 5'h2 == csrs_8_Index ? tlb_2_E : _GEN_291;
  wire  _GEN_293 = 5'h3 == csrs_8_Index ? tlb_3_E : _GEN_292;
  wire  _GEN_294 = 5'h4 == csrs_8_Index ? tlb_4_E : _GEN_293;
  wire  _GEN_295 = 5'h5 == csrs_8_Index ? tlb_5_E : _GEN_294;
  wire  _GEN_296 = 5'h6 == csrs_8_Index ? tlb_6_E : _GEN_295;
  wire  _GEN_297 = 5'h7 == csrs_8_Index ? tlb_7_E : _GEN_296;
  wire  _GEN_298 = 5'h8 == csrs_8_Index ? tlb_8_E : _GEN_297;
  wire  _GEN_299 = 5'h9 == csrs_8_Index ? tlb_9_E : _GEN_298;
  wire  _GEN_300 = 5'ha == csrs_8_Index ? tlb_10_E : _GEN_299;
  wire  _GEN_301 = 5'hb == csrs_8_Index ? tlb_11_E : _GEN_300;
  wire  _GEN_302 = 5'hc == csrs_8_Index ? tlb_12_E : _GEN_301;
  wire  _GEN_303 = 5'hd == csrs_8_Index ? tlb_13_E : _GEN_302;
  wire  _GEN_304 = 5'he == csrs_8_Index ? tlb_14_E : _GEN_303;
  wire  _GEN_305 = 5'hf == csrs_8_Index ? tlb_15_E : _GEN_304;
  wire  _GEN_306 = 5'h10 == csrs_8_Index ? tlb_16_E : _GEN_305;
  wire  _GEN_307 = 5'h11 == csrs_8_Index ? tlb_17_E : _GEN_306;
  wire  _GEN_308 = 5'h12 == csrs_8_Index ? tlb_18_E : _GEN_307;
  wire  _GEN_309 = 5'h13 == csrs_8_Index ? tlb_19_E : _GEN_308;
  wire  _GEN_310 = 5'h14 == csrs_8_Index ? tlb_20_E : _GEN_309;
  wire  _GEN_311 = 5'h15 == csrs_8_Index ? tlb_21_E : _GEN_310;
  wire  _GEN_312 = 5'h16 == csrs_8_Index ? tlb_22_E : _GEN_311;
  wire  _GEN_313 = 5'h17 == csrs_8_Index ? tlb_23_E : _GEN_312;
  wire  _GEN_314 = 5'h18 == csrs_8_Index ? tlb_24_E : _GEN_313;
  wire  _GEN_315 = 5'h19 == csrs_8_Index ? tlb_25_E : _GEN_314;
  wire  _GEN_316 = 5'h1a == csrs_8_Index ? tlb_26_E : _GEN_315;
  wire  _GEN_317 = 5'h1b == csrs_8_Index ? tlb_27_E : _GEN_316;
  wire  _GEN_318 = 5'h1c == csrs_8_Index ? tlb_28_E : _GEN_317;
  wire  _GEN_319 = 5'h1d == csrs_8_Index ? tlb_29_E : _GEN_318;
  wire  _GEN_320 = 5'h1e == csrs_8_Index ? tlb_30_E : _GEN_319;
  wire  _GEN_321 = 5'h1f == csrs_8_Index ? tlb_31_E : _GEN_320;
  wire [5:0] _GEN_323 = 5'h1 == csrs_8_Index ? tlb_1_PS : tlb_0_PS;
  wire [5:0] _GEN_324 = 5'h2 == csrs_8_Index ? tlb_2_PS : _GEN_323;
  wire [5:0] _GEN_325 = 5'h3 == csrs_8_Index ? tlb_3_PS : _GEN_324;
  wire [5:0] _GEN_326 = 5'h4 == csrs_8_Index ? tlb_4_PS : _GEN_325;
  wire [5:0] _GEN_327 = 5'h5 == csrs_8_Index ? tlb_5_PS : _GEN_326;
  wire [5:0] _GEN_328 = 5'h6 == csrs_8_Index ? tlb_6_PS : _GEN_327;
  wire [5:0] _GEN_329 = 5'h7 == csrs_8_Index ? tlb_7_PS : _GEN_328;
  wire [5:0] _GEN_330 = 5'h8 == csrs_8_Index ? tlb_8_PS : _GEN_329;
  wire [5:0] _GEN_331 = 5'h9 == csrs_8_Index ? tlb_9_PS : _GEN_330;
  wire [5:0] _GEN_332 = 5'ha == csrs_8_Index ? tlb_10_PS : _GEN_331;
  wire [5:0] _GEN_333 = 5'hb == csrs_8_Index ? tlb_11_PS : _GEN_332;
  wire [5:0] _GEN_334 = 5'hc == csrs_8_Index ? tlb_12_PS : _GEN_333;
  wire [5:0] _GEN_335 = 5'hd == csrs_8_Index ? tlb_13_PS : _GEN_334;
  wire [5:0] _GEN_336 = 5'he == csrs_8_Index ? tlb_14_PS : _GEN_335;
  wire [5:0] _GEN_337 = 5'hf == csrs_8_Index ? tlb_15_PS : _GEN_336;
  wire [5:0] _GEN_338 = 5'h10 == csrs_8_Index ? tlb_16_PS : _GEN_337;
  wire [5:0] _GEN_339 = 5'h11 == csrs_8_Index ? tlb_17_PS : _GEN_338;
  wire [5:0] _GEN_340 = 5'h12 == csrs_8_Index ? tlb_18_PS : _GEN_339;
  wire [5:0] _GEN_341 = 5'h13 == csrs_8_Index ? tlb_19_PS : _GEN_340;
  wire [5:0] _GEN_342 = 5'h14 == csrs_8_Index ? tlb_20_PS : _GEN_341;
  wire [5:0] _GEN_343 = 5'h15 == csrs_8_Index ? tlb_21_PS : _GEN_342;
  wire [5:0] _GEN_344 = 5'h16 == csrs_8_Index ? tlb_22_PS : _GEN_343;
  wire [5:0] _GEN_345 = 5'h17 == csrs_8_Index ? tlb_23_PS : _GEN_344;
  wire [5:0] _GEN_346 = 5'h18 == csrs_8_Index ? tlb_24_PS : _GEN_345;
  wire [5:0] _GEN_347 = 5'h19 == csrs_8_Index ? tlb_25_PS : _GEN_346;
  wire [5:0] _GEN_348 = 5'h1a == csrs_8_Index ? tlb_26_PS : _GEN_347;
  wire [5:0] _GEN_349 = 5'h1b == csrs_8_Index ? tlb_27_PS : _GEN_348;
  wire [5:0] _GEN_350 = 5'h1c == csrs_8_Index ? tlb_28_PS : _GEN_349;
  wire [5:0] _GEN_351 = 5'h1d == csrs_8_Index ? tlb_29_PS : _GEN_350;
  wire [5:0] _GEN_352 = 5'h1e == csrs_8_Index ? tlb_30_PS : _GEN_351;
  wire [5:0] _GEN_353 = 5'h1f == csrs_8_Index ? tlb_31_PS : _GEN_352;
  wire [18:0] _GEN_355 = 5'h1 == csrs_8_Index ? tlb_1_VPPN : tlb_0_VPPN;
  wire [18:0] _GEN_356 = 5'h2 == csrs_8_Index ? tlb_2_VPPN : _GEN_355;
  wire [18:0] _GEN_357 = 5'h3 == csrs_8_Index ? tlb_3_VPPN : _GEN_356;
  wire [18:0] _GEN_358 = 5'h4 == csrs_8_Index ? tlb_4_VPPN : _GEN_357;
  wire [18:0] _GEN_359 = 5'h5 == csrs_8_Index ? tlb_5_VPPN : _GEN_358;
  wire [18:0] _GEN_360 = 5'h6 == csrs_8_Index ? tlb_6_VPPN : _GEN_359;
  wire [18:0] _GEN_361 = 5'h7 == csrs_8_Index ? tlb_7_VPPN : _GEN_360;
  wire [18:0] _GEN_362 = 5'h8 == csrs_8_Index ? tlb_8_VPPN : _GEN_361;
  wire [18:0] _GEN_363 = 5'h9 == csrs_8_Index ? tlb_9_VPPN : _GEN_362;
  wire [18:0] _GEN_364 = 5'ha == csrs_8_Index ? tlb_10_VPPN : _GEN_363;
  wire [18:0] _GEN_365 = 5'hb == csrs_8_Index ? tlb_11_VPPN : _GEN_364;
  wire [18:0] _GEN_366 = 5'hc == csrs_8_Index ? tlb_12_VPPN : _GEN_365;
  wire [18:0] _GEN_367 = 5'hd == csrs_8_Index ? tlb_13_VPPN : _GEN_366;
  wire [18:0] _GEN_368 = 5'he == csrs_8_Index ? tlb_14_VPPN : _GEN_367;
  wire [18:0] _GEN_369 = 5'hf == csrs_8_Index ? tlb_15_VPPN : _GEN_368;
  wire [18:0] _GEN_370 = 5'h10 == csrs_8_Index ? tlb_16_VPPN : _GEN_369;
  wire [18:0] _GEN_371 = 5'h11 == csrs_8_Index ? tlb_17_VPPN : _GEN_370;
  wire [18:0] _GEN_372 = 5'h12 == csrs_8_Index ? tlb_18_VPPN : _GEN_371;
  wire [18:0] _GEN_373 = 5'h13 == csrs_8_Index ? tlb_19_VPPN : _GEN_372;
  wire [18:0] _GEN_374 = 5'h14 == csrs_8_Index ? tlb_20_VPPN : _GEN_373;
  wire [18:0] _GEN_375 = 5'h15 == csrs_8_Index ? tlb_21_VPPN : _GEN_374;
  wire [18:0] _GEN_376 = 5'h16 == csrs_8_Index ? tlb_22_VPPN : _GEN_375;
  wire [18:0] _GEN_377 = 5'h17 == csrs_8_Index ? tlb_23_VPPN : _GEN_376;
  wire [18:0] _GEN_378 = 5'h18 == csrs_8_Index ? tlb_24_VPPN : _GEN_377;
  wire [18:0] _GEN_379 = 5'h19 == csrs_8_Index ? tlb_25_VPPN : _GEN_378;
  wire [18:0] _GEN_380 = 5'h1a == csrs_8_Index ? tlb_26_VPPN : _GEN_379;
  wire [18:0] _GEN_381 = 5'h1b == csrs_8_Index ? tlb_27_VPPN : _GEN_380;
  wire [18:0] _GEN_382 = 5'h1c == csrs_8_Index ? tlb_28_VPPN : _GEN_381;
  wire [18:0] _GEN_383 = 5'h1d == csrs_8_Index ? tlb_29_VPPN : _GEN_382;
  wire [18:0] _GEN_384 = 5'h1e == csrs_8_Index ? tlb_30_VPPN : _GEN_383;
  wire [18:0] _GEN_385 = 5'h1f == csrs_8_Index ? tlb_31_VPPN : _GEN_384;
  wire [19:0] _GEN_387 = 5'h1 == csrs_8_Index ? tlb_1_P0_PPN : tlb_0_P0_PPN;
  wire [19:0] _GEN_388 = 5'h2 == csrs_8_Index ? tlb_2_P0_PPN : _GEN_387;
  wire [19:0] _GEN_389 = 5'h3 == csrs_8_Index ? tlb_3_P0_PPN : _GEN_388;
  wire [19:0] _GEN_390 = 5'h4 == csrs_8_Index ? tlb_4_P0_PPN : _GEN_389;
  wire [19:0] _GEN_391 = 5'h5 == csrs_8_Index ? tlb_5_P0_PPN : _GEN_390;
  wire [19:0] _GEN_392 = 5'h6 == csrs_8_Index ? tlb_6_P0_PPN : _GEN_391;
  wire [19:0] _GEN_393 = 5'h7 == csrs_8_Index ? tlb_7_P0_PPN : _GEN_392;
  wire [19:0] _GEN_394 = 5'h8 == csrs_8_Index ? tlb_8_P0_PPN : _GEN_393;
  wire [19:0] _GEN_395 = 5'h9 == csrs_8_Index ? tlb_9_P0_PPN : _GEN_394;
  wire [19:0] _GEN_396 = 5'ha == csrs_8_Index ? tlb_10_P0_PPN : _GEN_395;
  wire [19:0] _GEN_397 = 5'hb == csrs_8_Index ? tlb_11_P0_PPN : _GEN_396;
  wire [19:0] _GEN_398 = 5'hc == csrs_8_Index ? tlb_12_P0_PPN : _GEN_397;
  wire [19:0] _GEN_399 = 5'hd == csrs_8_Index ? tlb_13_P0_PPN : _GEN_398;
  wire [19:0] _GEN_400 = 5'he == csrs_8_Index ? tlb_14_P0_PPN : _GEN_399;
  wire [19:0] _GEN_401 = 5'hf == csrs_8_Index ? tlb_15_P0_PPN : _GEN_400;
  wire [19:0] _GEN_402 = 5'h10 == csrs_8_Index ? tlb_16_P0_PPN : _GEN_401;
  wire [19:0] _GEN_403 = 5'h11 == csrs_8_Index ? tlb_17_P0_PPN : _GEN_402;
  wire [19:0] _GEN_404 = 5'h12 == csrs_8_Index ? tlb_18_P0_PPN : _GEN_403;
  wire [19:0] _GEN_405 = 5'h13 == csrs_8_Index ? tlb_19_P0_PPN : _GEN_404;
  wire [19:0] _GEN_406 = 5'h14 == csrs_8_Index ? tlb_20_P0_PPN : _GEN_405;
  wire [19:0] _GEN_407 = 5'h15 == csrs_8_Index ? tlb_21_P0_PPN : _GEN_406;
  wire [19:0] _GEN_408 = 5'h16 == csrs_8_Index ? tlb_22_P0_PPN : _GEN_407;
  wire [19:0] _GEN_409 = 5'h17 == csrs_8_Index ? tlb_23_P0_PPN : _GEN_408;
  wire [19:0] _GEN_410 = 5'h18 == csrs_8_Index ? tlb_24_P0_PPN : _GEN_409;
  wire [19:0] _GEN_411 = 5'h19 == csrs_8_Index ? tlb_25_P0_PPN : _GEN_410;
  wire [19:0] _GEN_412 = 5'h1a == csrs_8_Index ? tlb_26_P0_PPN : _GEN_411;
  wire [19:0] _GEN_413 = 5'h1b == csrs_8_Index ? tlb_27_P0_PPN : _GEN_412;
  wire [19:0] _GEN_414 = 5'h1c == csrs_8_Index ? tlb_28_P0_PPN : _GEN_413;
  wire [19:0] _GEN_415 = 5'h1d == csrs_8_Index ? tlb_29_P0_PPN : _GEN_414;
  wire [19:0] _GEN_416 = 5'h1e == csrs_8_Index ? tlb_30_P0_PPN : _GEN_415;
  wire [19:0] _GEN_417 = 5'h1f == csrs_8_Index ? tlb_31_P0_PPN : _GEN_416;
  wire  _GEN_419 = 5'h1 == csrs_8_Index ? tlb_1_G : tlb_0_G;
  wire  _GEN_420 = 5'h2 == csrs_8_Index ? tlb_2_G : _GEN_419;
  wire  _GEN_421 = 5'h3 == csrs_8_Index ? tlb_3_G : _GEN_420;
  wire  _GEN_422 = 5'h4 == csrs_8_Index ? tlb_4_G : _GEN_421;
  wire  _GEN_423 = 5'h5 == csrs_8_Index ? tlb_5_G : _GEN_422;
  wire  _GEN_424 = 5'h6 == csrs_8_Index ? tlb_6_G : _GEN_423;
  wire  _GEN_425 = 5'h7 == csrs_8_Index ? tlb_7_G : _GEN_424;
  wire  _GEN_426 = 5'h8 == csrs_8_Index ? tlb_8_G : _GEN_425;
  wire  _GEN_427 = 5'h9 == csrs_8_Index ? tlb_9_G : _GEN_426;
  wire  _GEN_428 = 5'ha == csrs_8_Index ? tlb_10_G : _GEN_427;
  wire  _GEN_429 = 5'hb == csrs_8_Index ? tlb_11_G : _GEN_428;
  wire  _GEN_430 = 5'hc == csrs_8_Index ? tlb_12_G : _GEN_429;
  wire  _GEN_431 = 5'hd == csrs_8_Index ? tlb_13_G : _GEN_430;
  wire  _GEN_432 = 5'he == csrs_8_Index ? tlb_14_G : _GEN_431;
  wire  _GEN_433 = 5'hf == csrs_8_Index ? tlb_15_G : _GEN_432;
  wire  _GEN_434 = 5'h10 == csrs_8_Index ? tlb_16_G : _GEN_433;
  wire  _GEN_435 = 5'h11 == csrs_8_Index ? tlb_17_G : _GEN_434;
  wire  _GEN_436 = 5'h12 == csrs_8_Index ? tlb_18_G : _GEN_435;
  wire  _GEN_437 = 5'h13 == csrs_8_Index ? tlb_19_G : _GEN_436;
  wire  _GEN_438 = 5'h14 == csrs_8_Index ? tlb_20_G : _GEN_437;
  wire  _GEN_439 = 5'h15 == csrs_8_Index ? tlb_21_G : _GEN_438;
  wire  _GEN_440 = 5'h16 == csrs_8_Index ? tlb_22_G : _GEN_439;
  wire  _GEN_441 = 5'h17 == csrs_8_Index ? tlb_23_G : _GEN_440;
  wire  _GEN_442 = 5'h18 == csrs_8_Index ? tlb_24_G : _GEN_441;
  wire  _GEN_443 = 5'h19 == csrs_8_Index ? tlb_25_G : _GEN_442;
  wire  _GEN_444 = 5'h1a == csrs_8_Index ? tlb_26_G : _GEN_443;
  wire  _GEN_445 = 5'h1b == csrs_8_Index ? tlb_27_G : _GEN_444;
  wire  _GEN_446 = 5'h1c == csrs_8_Index ? tlb_28_G : _GEN_445;
  wire  _GEN_447 = 5'h1d == csrs_8_Index ? tlb_29_G : _GEN_446;
  wire  _GEN_448 = 5'h1e == csrs_8_Index ? tlb_30_G : _GEN_447;
  wire  _GEN_449 = 5'h1f == csrs_8_Index ? tlb_31_G : _GEN_448;
  wire [1:0] _GEN_451 = 5'h1 == csrs_8_Index ? tlb_1_P0_MAT : tlb_0_P0_MAT;
  wire [1:0] _GEN_452 = 5'h2 == csrs_8_Index ? tlb_2_P0_MAT : _GEN_451;
  wire [1:0] _GEN_453 = 5'h3 == csrs_8_Index ? tlb_3_P0_MAT : _GEN_452;
  wire [1:0] _GEN_454 = 5'h4 == csrs_8_Index ? tlb_4_P0_MAT : _GEN_453;
  wire [1:0] _GEN_455 = 5'h5 == csrs_8_Index ? tlb_5_P0_MAT : _GEN_454;
  wire [1:0] _GEN_456 = 5'h6 == csrs_8_Index ? tlb_6_P0_MAT : _GEN_455;
  wire [1:0] _GEN_457 = 5'h7 == csrs_8_Index ? tlb_7_P0_MAT : _GEN_456;
  wire [1:0] _GEN_458 = 5'h8 == csrs_8_Index ? tlb_8_P0_MAT : _GEN_457;
  wire [1:0] _GEN_459 = 5'h9 == csrs_8_Index ? tlb_9_P0_MAT : _GEN_458;
  wire [1:0] _GEN_460 = 5'ha == csrs_8_Index ? tlb_10_P0_MAT : _GEN_459;
  wire [1:0] _GEN_461 = 5'hb == csrs_8_Index ? tlb_11_P0_MAT : _GEN_460;
  wire [1:0] _GEN_462 = 5'hc == csrs_8_Index ? tlb_12_P0_MAT : _GEN_461;
  wire [1:0] _GEN_463 = 5'hd == csrs_8_Index ? tlb_13_P0_MAT : _GEN_462;
  wire [1:0] _GEN_464 = 5'he == csrs_8_Index ? tlb_14_P0_MAT : _GEN_463;
  wire [1:0] _GEN_465 = 5'hf == csrs_8_Index ? tlb_15_P0_MAT : _GEN_464;
  wire [1:0] _GEN_466 = 5'h10 == csrs_8_Index ? tlb_16_P0_MAT : _GEN_465;
  wire [1:0] _GEN_467 = 5'h11 == csrs_8_Index ? tlb_17_P0_MAT : _GEN_466;
  wire [1:0] _GEN_468 = 5'h12 == csrs_8_Index ? tlb_18_P0_MAT : _GEN_467;
  wire [1:0] _GEN_469 = 5'h13 == csrs_8_Index ? tlb_19_P0_MAT : _GEN_468;
  wire [1:0] _GEN_470 = 5'h14 == csrs_8_Index ? tlb_20_P0_MAT : _GEN_469;
  wire [1:0] _GEN_471 = 5'h15 == csrs_8_Index ? tlb_21_P0_MAT : _GEN_470;
  wire [1:0] _GEN_472 = 5'h16 == csrs_8_Index ? tlb_22_P0_MAT : _GEN_471;
  wire [1:0] _GEN_473 = 5'h17 == csrs_8_Index ? tlb_23_P0_MAT : _GEN_472;
  wire [1:0] _GEN_474 = 5'h18 == csrs_8_Index ? tlb_24_P0_MAT : _GEN_473;
  wire [1:0] _GEN_475 = 5'h19 == csrs_8_Index ? tlb_25_P0_MAT : _GEN_474;
  wire [1:0] _GEN_476 = 5'h1a == csrs_8_Index ? tlb_26_P0_MAT : _GEN_475;
  wire [1:0] _GEN_477 = 5'h1b == csrs_8_Index ? tlb_27_P0_MAT : _GEN_476;
  wire [1:0] _GEN_478 = 5'h1c == csrs_8_Index ? tlb_28_P0_MAT : _GEN_477;
  wire [1:0] _GEN_479 = 5'h1d == csrs_8_Index ? tlb_29_P0_MAT : _GEN_478;
  wire [1:0] _GEN_480 = 5'h1e == csrs_8_Index ? tlb_30_P0_MAT : _GEN_479;
  wire [1:0] _GEN_481 = 5'h1f == csrs_8_Index ? tlb_31_P0_MAT : _GEN_480;
  wire [1:0] _GEN_483 = 5'h1 == csrs_8_Index ? tlb_1_P0_PLV : tlb_0_P0_PLV;
  wire [1:0] _GEN_484 = 5'h2 == csrs_8_Index ? tlb_2_P0_PLV : _GEN_483;
  wire [1:0] _GEN_485 = 5'h3 == csrs_8_Index ? tlb_3_P0_PLV : _GEN_484;
  wire [1:0] _GEN_486 = 5'h4 == csrs_8_Index ? tlb_4_P0_PLV : _GEN_485;
  wire [1:0] _GEN_487 = 5'h5 == csrs_8_Index ? tlb_5_P0_PLV : _GEN_486;
  wire [1:0] _GEN_488 = 5'h6 == csrs_8_Index ? tlb_6_P0_PLV : _GEN_487;
  wire [1:0] _GEN_489 = 5'h7 == csrs_8_Index ? tlb_7_P0_PLV : _GEN_488;
  wire [1:0] _GEN_490 = 5'h8 == csrs_8_Index ? tlb_8_P0_PLV : _GEN_489;
  wire [1:0] _GEN_491 = 5'h9 == csrs_8_Index ? tlb_9_P0_PLV : _GEN_490;
  wire [1:0] _GEN_492 = 5'ha == csrs_8_Index ? tlb_10_P0_PLV : _GEN_491;
  wire [1:0] _GEN_493 = 5'hb == csrs_8_Index ? tlb_11_P0_PLV : _GEN_492;
  wire [1:0] _GEN_494 = 5'hc == csrs_8_Index ? tlb_12_P0_PLV : _GEN_493;
  wire [1:0] _GEN_495 = 5'hd == csrs_8_Index ? tlb_13_P0_PLV : _GEN_494;
  wire [1:0] _GEN_496 = 5'he == csrs_8_Index ? tlb_14_P0_PLV : _GEN_495;
  wire [1:0] _GEN_497 = 5'hf == csrs_8_Index ? tlb_15_P0_PLV : _GEN_496;
  wire [1:0] _GEN_498 = 5'h10 == csrs_8_Index ? tlb_16_P0_PLV : _GEN_497;
  wire [1:0] _GEN_499 = 5'h11 == csrs_8_Index ? tlb_17_P0_PLV : _GEN_498;
  wire [1:0] _GEN_500 = 5'h12 == csrs_8_Index ? tlb_18_P0_PLV : _GEN_499;
  wire [1:0] _GEN_501 = 5'h13 == csrs_8_Index ? tlb_19_P0_PLV : _GEN_500;
  wire [1:0] _GEN_502 = 5'h14 == csrs_8_Index ? tlb_20_P0_PLV : _GEN_501;
  wire [1:0] _GEN_503 = 5'h15 == csrs_8_Index ? tlb_21_P0_PLV : _GEN_502;
  wire [1:0] _GEN_504 = 5'h16 == csrs_8_Index ? tlb_22_P0_PLV : _GEN_503;
  wire [1:0] _GEN_505 = 5'h17 == csrs_8_Index ? tlb_23_P0_PLV : _GEN_504;
  wire [1:0] _GEN_506 = 5'h18 == csrs_8_Index ? tlb_24_P0_PLV : _GEN_505;
  wire [1:0] _GEN_507 = 5'h19 == csrs_8_Index ? tlb_25_P0_PLV : _GEN_506;
  wire [1:0] _GEN_508 = 5'h1a == csrs_8_Index ? tlb_26_P0_PLV : _GEN_507;
  wire [1:0] _GEN_509 = 5'h1b == csrs_8_Index ? tlb_27_P0_PLV : _GEN_508;
  wire [1:0] _GEN_510 = 5'h1c == csrs_8_Index ? tlb_28_P0_PLV : _GEN_509;
  wire [1:0] _GEN_511 = 5'h1d == csrs_8_Index ? tlb_29_P0_PLV : _GEN_510;
  wire [1:0] _GEN_512 = 5'h1e == csrs_8_Index ? tlb_30_P0_PLV : _GEN_511;
  wire [1:0] _GEN_513 = 5'h1f == csrs_8_Index ? tlb_31_P0_PLV : _GEN_512;
  wire  _GEN_515 = 5'h1 == csrs_8_Index ? tlb_1_P0_D : tlb_0_P0_D;
  wire  _GEN_516 = 5'h2 == csrs_8_Index ? tlb_2_P0_D : _GEN_515;
  wire  _GEN_517 = 5'h3 == csrs_8_Index ? tlb_3_P0_D : _GEN_516;
  wire  _GEN_518 = 5'h4 == csrs_8_Index ? tlb_4_P0_D : _GEN_517;
  wire  _GEN_519 = 5'h5 == csrs_8_Index ? tlb_5_P0_D : _GEN_518;
  wire  _GEN_520 = 5'h6 == csrs_8_Index ? tlb_6_P0_D : _GEN_519;
  wire  _GEN_521 = 5'h7 == csrs_8_Index ? tlb_7_P0_D : _GEN_520;
  wire  _GEN_522 = 5'h8 == csrs_8_Index ? tlb_8_P0_D : _GEN_521;
  wire  _GEN_523 = 5'h9 == csrs_8_Index ? tlb_9_P0_D : _GEN_522;
  wire  _GEN_524 = 5'ha == csrs_8_Index ? tlb_10_P0_D : _GEN_523;
  wire  _GEN_525 = 5'hb == csrs_8_Index ? tlb_11_P0_D : _GEN_524;
  wire  _GEN_526 = 5'hc == csrs_8_Index ? tlb_12_P0_D : _GEN_525;
  wire  _GEN_527 = 5'hd == csrs_8_Index ? tlb_13_P0_D : _GEN_526;
  wire  _GEN_528 = 5'he == csrs_8_Index ? tlb_14_P0_D : _GEN_527;
  wire  _GEN_529 = 5'hf == csrs_8_Index ? tlb_15_P0_D : _GEN_528;
  wire  _GEN_530 = 5'h10 == csrs_8_Index ? tlb_16_P0_D : _GEN_529;
  wire  _GEN_531 = 5'h11 == csrs_8_Index ? tlb_17_P0_D : _GEN_530;
  wire  _GEN_532 = 5'h12 == csrs_8_Index ? tlb_18_P0_D : _GEN_531;
  wire  _GEN_533 = 5'h13 == csrs_8_Index ? tlb_19_P0_D : _GEN_532;
  wire  _GEN_534 = 5'h14 == csrs_8_Index ? tlb_20_P0_D : _GEN_533;
  wire  _GEN_535 = 5'h15 == csrs_8_Index ? tlb_21_P0_D : _GEN_534;
  wire  _GEN_536 = 5'h16 == csrs_8_Index ? tlb_22_P0_D : _GEN_535;
  wire  _GEN_537 = 5'h17 == csrs_8_Index ? tlb_23_P0_D : _GEN_536;
  wire  _GEN_538 = 5'h18 == csrs_8_Index ? tlb_24_P0_D : _GEN_537;
  wire  _GEN_539 = 5'h19 == csrs_8_Index ? tlb_25_P0_D : _GEN_538;
  wire  _GEN_540 = 5'h1a == csrs_8_Index ? tlb_26_P0_D : _GEN_539;
  wire  _GEN_541 = 5'h1b == csrs_8_Index ? tlb_27_P0_D : _GEN_540;
  wire  _GEN_542 = 5'h1c == csrs_8_Index ? tlb_28_P0_D : _GEN_541;
  wire  _GEN_543 = 5'h1d == csrs_8_Index ? tlb_29_P0_D : _GEN_542;
  wire  _GEN_544 = 5'h1e == csrs_8_Index ? tlb_30_P0_D : _GEN_543;
  wire  _GEN_545 = 5'h1f == csrs_8_Index ? tlb_31_P0_D : _GEN_544;
  wire  _GEN_547 = 5'h1 == csrs_8_Index ? tlb_1_P0_V : tlb_0_P0_V;
  wire  _GEN_548 = 5'h2 == csrs_8_Index ? tlb_2_P0_V : _GEN_547;
  wire  _GEN_549 = 5'h3 == csrs_8_Index ? tlb_3_P0_V : _GEN_548;
  wire  _GEN_550 = 5'h4 == csrs_8_Index ? tlb_4_P0_V : _GEN_549;
  wire  _GEN_551 = 5'h5 == csrs_8_Index ? tlb_5_P0_V : _GEN_550;
  wire  _GEN_552 = 5'h6 == csrs_8_Index ? tlb_6_P0_V : _GEN_551;
  wire  _GEN_553 = 5'h7 == csrs_8_Index ? tlb_7_P0_V : _GEN_552;
  wire  _GEN_554 = 5'h8 == csrs_8_Index ? tlb_8_P0_V : _GEN_553;
  wire  _GEN_555 = 5'h9 == csrs_8_Index ? tlb_9_P0_V : _GEN_554;
  wire  _GEN_556 = 5'ha == csrs_8_Index ? tlb_10_P0_V : _GEN_555;
  wire  _GEN_557 = 5'hb == csrs_8_Index ? tlb_11_P0_V : _GEN_556;
  wire  _GEN_558 = 5'hc == csrs_8_Index ? tlb_12_P0_V : _GEN_557;
  wire  _GEN_559 = 5'hd == csrs_8_Index ? tlb_13_P0_V : _GEN_558;
  wire  _GEN_560 = 5'he == csrs_8_Index ? tlb_14_P0_V : _GEN_559;
  wire  _GEN_561 = 5'hf == csrs_8_Index ? tlb_15_P0_V : _GEN_560;
  wire  _GEN_562 = 5'h10 == csrs_8_Index ? tlb_16_P0_V : _GEN_561;
  wire  _GEN_563 = 5'h11 == csrs_8_Index ? tlb_17_P0_V : _GEN_562;
  wire  _GEN_564 = 5'h12 == csrs_8_Index ? tlb_18_P0_V : _GEN_563;
  wire  _GEN_565 = 5'h13 == csrs_8_Index ? tlb_19_P0_V : _GEN_564;
  wire  _GEN_566 = 5'h14 == csrs_8_Index ? tlb_20_P0_V : _GEN_565;
  wire  _GEN_567 = 5'h15 == csrs_8_Index ? tlb_21_P0_V : _GEN_566;
  wire  _GEN_568 = 5'h16 == csrs_8_Index ? tlb_22_P0_V : _GEN_567;
  wire  _GEN_569 = 5'h17 == csrs_8_Index ? tlb_23_P0_V : _GEN_568;
  wire  _GEN_570 = 5'h18 == csrs_8_Index ? tlb_24_P0_V : _GEN_569;
  wire  _GEN_571 = 5'h19 == csrs_8_Index ? tlb_25_P0_V : _GEN_570;
  wire  _GEN_572 = 5'h1a == csrs_8_Index ? tlb_26_P0_V : _GEN_571;
  wire  _GEN_573 = 5'h1b == csrs_8_Index ? tlb_27_P0_V : _GEN_572;
  wire  _GEN_574 = 5'h1c == csrs_8_Index ? tlb_28_P0_V : _GEN_573;
  wire  _GEN_575 = 5'h1d == csrs_8_Index ? tlb_29_P0_V : _GEN_574;
  wire  _GEN_576 = 5'h1e == csrs_8_Index ? tlb_30_P0_V : _GEN_575;
  wire  _GEN_577 = 5'h1f == csrs_8_Index ? tlb_31_P0_V : _GEN_576;
  wire [19:0] _GEN_579 = 5'h1 == csrs_8_Index ? tlb_1_P1_PPN : tlb_0_P1_PPN;
  wire [19:0] _GEN_580 = 5'h2 == csrs_8_Index ? tlb_2_P1_PPN : _GEN_579;
  wire [19:0] _GEN_581 = 5'h3 == csrs_8_Index ? tlb_3_P1_PPN : _GEN_580;
  wire [19:0] _GEN_582 = 5'h4 == csrs_8_Index ? tlb_4_P1_PPN : _GEN_581;
  wire [19:0] _GEN_583 = 5'h5 == csrs_8_Index ? tlb_5_P1_PPN : _GEN_582;
  wire [19:0] _GEN_584 = 5'h6 == csrs_8_Index ? tlb_6_P1_PPN : _GEN_583;
  wire [19:0] _GEN_585 = 5'h7 == csrs_8_Index ? tlb_7_P1_PPN : _GEN_584;
  wire [19:0] _GEN_586 = 5'h8 == csrs_8_Index ? tlb_8_P1_PPN : _GEN_585;
  wire [19:0] _GEN_587 = 5'h9 == csrs_8_Index ? tlb_9_P1_PPN : _GEN_586;
  wire [19:0] _GEN_588 = 5'ha == csrs_8_Index ? tlb_10_P1_PPN : _GEN_587;
  wire [19:0] _GEN_589 = 5'hb == csrs_8_Index ? tlb_11_P1_PPN : _GEN_588;
  wire [19:0] _GEN_590 = 5'hc == csrs_8_Index ? tlb_12_P1_PPN : _GEN_589;
  wire [19:0] _GEN_591 = 5'hd == csrs_8_Index ? tlb_13_P1_PPN : _GEN_590;
  wire [19:0] _GEN_592 = 5'he == csrs_8_Index ? tlb_14_P1_PPN : _GEN_591;
  wire [19:0] _GEN_593 = 5'hf == csrs_8_Index ? tlb_15_P1_PPN : _GEN_592;
  wire [19:0] _GEN_594 = 5'h10 == csrs_8_Index ? tlb_16_P1_PPN : _GEN_593;
  wire [19:0] _GEN_595 = 5'h11 == csrs_8_Index ? tlb_17_P1_PPN : _GEN_594;
  wire [19:0] _GEN_596 = 5'h12 == csrs_8_Index ? tlb_18_P1_PPN : _GEN_595;
  wire [19:0] _GEN_597 = 5'h13 == csrs_8_Index ? tlb_19_P1_PPN : _GEN_596;
  wire [19:0] _GEN_598 = 5'h14 == csrs_8_Index ? tlb_20_P1_PPN : _GEN_597;
  wire [19:0] _GEN_599 = 5'h15 == csrs_8_Index ? tlb_21_P1_PPN : _GEN_598;
  wire [19:0] _GEN_600 = 5'h16 == csrs_8_Index ? tlb_22_P1_PPN : _GEN_599;
  wire [19:0] _GEN_601 = 5'h17 == csrs_8_Index ? tlb_23_P1_PPN : _GEN_600;
  wire [19:0] _GEN_602 = 5'h18 == csrs_8_Index ? tlb_24_P1_PPN : _GEN_601;
  wire [19:0] _GEN_603 = 5'h19 == csrs_8_Index ? tlb_25_P1_PPN : _GEN_602;
  wire [19:0] _GEN_604 = 5'h1a == csrs_8_Index ? tlb_26_P1_PPN : _GEN_603;
  wire [19:0] _GEN_605 = 5'h1b == csrs_8_Index ? tlb_27_P1_PPN : _GEN_604;
  wire [19:0] _GEN_606 = 5'h1c == csrs_8_Index ? tlb_28_P1_PPN : _GEN_605;
  wire [19:0] _GEN_607 = 5'h1d == csrs_8_Index ? tlb_29_P1_PPN : _GEN_606;
  wire [19:0] _GEN_608 = 5'h1e == csrs_8_Index ? tlb_30_P1_PPN : _GEN_607;
  wire [19:0] _GEN_609 = 5'h1f == csrs_8_Index ? tlb_31_P1_PPN : _GEN_608;
  wire [1:0] _GEN_611 = 5'h1 == csrs_8_Index ? tlb_1_P1_MAT : tlb_0_P1_MAT;
  wire [1:0] _GEN_612 = 5'h2 == csrs_8_Index ? tlb_2_P1_MAT : _GEN_611;
  wire [1:0] _GEN_613 = 5'h3 == csrs_8_Index ? tlb_3_P1_MAT : _GEN_612;
  wire [1:0] _GEN_614 = 5'h4 == csrs_8_Index ? tlb_4_P1_MAT : _GEN_613;
  wire [1:0] _GEN_615 = 5'h5 == csrs_8_Index ? tlb_5_P1_MAT : _GEN_614;
  wire [1:0] _GEN_616 = 5'h6 == csrs_8_Index ? tlb_6_P1_MAT : _GEN_615;
  wire [1:0] _GEN_617 = 5'h7 == csrs_8_Index ? tlb_7_P1_MAT : _GEN_616;
  wire [1:0] _GEN_618 = 5'h8 == csrs_8_Index ? tlb_8_P1_MAT : _GEN_617;
  wire [1:0] _GEN_619 = 5'h9 == csrs_8_Index ? tlb_9_P1_MAT : _GEN_618;
  wire [1:0] _GEN_620 = 5'ha == csrs_8_Index ? tlb_10_P1_MAT : _GEN_619;
  wire [1:0] _GEN_621 = 5'hb == csrs_8_Index ? tlb_11_P1_MAT : _GEN_620;
  wire [1:0] _GEN_622 = 5'hc == csrs_8_Index ? tlb_12_P1_MAT : _GEN_621;
  wire [1:0] _GEN_623 = 5'hd == csrs_8_Index ? tlb_13_P1_MAT : _GEN_622;
  wire [1:0] _GEN_624 = 5'he == csrs_8_Index ? tlb_14_P1_MAT : _GEN_623;
  wire [1:0] _GEN_625 = 5'hf == csrs_8_Index ? tlb_15_P1_MAT : _GEN_624;
  wire [1:0] _GEN_626 = 5'h10 == csrs_8_Index ? tlb_16_P1_MAT : _GEN_625;
  wire [1:0] _GEN_627 = 5'h11 == csrs_8_Index ? tlb_17_P1_MAT : _GEN_626;
  wire [1:0] _GEN_628 = 5'h12 == csrs_8_Index ? tlb_18_P1_MAT : _GEN_627;
  wire [1:0] _GEN_629 = 5'h13 == csrs_8_Index ? tlb_19_P1_MAT : _GEN_628;
  wire [1:0] _GEN_630 = 5'h14 == csrs_8_Index ? tlb_20_P1_MAT : _GEN_629;
  wire [1:0] _GEN_631 = 5'h15 == csrs_8_Index ? tlb_21_P1_MAT : _GEN_630;
  wire [1:0] _GEN_632 = 5'h16 == csrs_8_Index ? tlb_22_P1_MAT : _GEN_631;
  wire [1:0] _GEN_633 = 5'h17 == csrs_8_Index ? tlb_23_P1_MAT : _GEN_632;
  wire [1:0] _GEN_634 = 5'h18 == csrs_8_Index ? tlb_24_P1_MAT : _GEN_633;
  wire [1:0] _GEN_635 = 5'h19 == csrs_8_Index ? tlb_25_P1_MAT : _GEN_634;
  wire [1:0] _GEN_636 = 5'h1a == csrs_8_Index ? tlb_26_P1_MAT : _GEN_635;
  wire [1:0] _GEN_637 = 5'h1b == csrs_8_Index ? tlb_27_P1_MAT : _GEN_636;
  wire [1:0] _GEN_638 = 5'h1c == csrs_8_Index ? tlb_28_P1_MAT : _GEN_637;
  wire [1:0] _GEN_639 = 5'h1d == csrs_8_Index ? tlb_29_P1_MAT : _GEN_638;
  wire [1:0] _GEN_640 = 5'h1e == csrs_8_Index ? tlb_30_P1_MAT : _GEN_639;
  wire [1:0] _GEN_641 = 5'h1f == csrs_8_Index ? tlb_31_P1_MAT : _GEN_640;
  wire [1:0] _GEN_643 = 5'h1 == csrs_8_Index ? tlb_1_P1_PLV : tlb_0_P1_PLV;
  wire [1:0] _GEN_644 = 5'h2 == csrs_8_Index ? tlb_2_P1_PLV : _GEN_643;
  wire [1:0] _GEN_645 = 5'h3 == csrs_8_Index ? tlb_3_P1_PLV : _GEN_644;
  wire [1:0] _GEN_646 = 5'h4 == csrs_8_Index ? tlb_4_P1_PLV : _GEN_645;
  wire [1:0] _GEN_647 = 5'h5 == csrs_8_Index ? tlb_5_P1_PLV : _GEN_646;
  wire [1:0] _GEN_648 = 5'h6 == csrs_8_Index ? tlb_6_P1_PLV : _GEN_647;
  wire [1:0] _GEN_649 = 5'h7 == csrs_8_Index ? tlb_7_P1_PLV : _GEN_648;
  wire [1:0] _GEN_650 = 5'h8 == csrs_8_Index ? tlb_8_P1_PLV : _GEN_649;
  wire [1:0] _GEN_651 = 5'h9 == csrs_8_Index ? tlb_9_P1_PLV : _GEN_650;
  wire [1:0] _GEN_652 = 5'ha == csrs_8_Index ? tlb_10_P1_PLV : _GEN_651;
  wire [1:0] _GEN_653 = 5'hb == csrs_8_Index ? tlb_11_P1_PLV : _GEN_652;
  wire [1:0] _GEN_654 = 5'hc == csrs_8_Index ? tlb_12_P1_PLV : _GEN_653;
  wire [1:0] _GEN_655 = 5'hd == csrs_8_Index ? tlb_13_P1_PLV : _GEN_654;
  wire [1:0] _GEN_656 = 5'he == csrs_8_Index ? tlb_14_P1_PLV : _GEN_655;
  wire [1:0] _GEN_657 = 5'hf == csrs_8_Index ? tlb_15_P1_PLV : _GEN_656;
  wire [1:0] _GEN_658 = 5'h10 == csrs_8_Index ? tlb_16_P1_PLV : _GEN_657;
  wire [1:0] _GEN_659 = 5'h11 == csrs_8_Index ? tlb_17_P1_PLV : _GEN_658;
  wire [1:0] _GEN_660 = 5'h12 == csrs_8_Index ? tlb_18_P1_PLV : _GEN_659;
  wire [1:0] _GEN_661 = 5'h13 == csrs_8_Index ? tlb_19_P1_PLV : _GEN_660;
  wire [1:0] _GEN_662 = 5'h14 == csrs_8_Index ? tlb_20_P1_PLV : _GEN_661;
  wire [1:0] _GEN_663 = 5'h15 == csrs_8_Index ? tlb_21_P1_PLV : _GEN_662;
  wire [1:0] _GEN_664 = 5'h16 == csrs_8_Index ? tlb_22_P1_PLV : _GEN_663;
  wire [1:0] _GEN_665 = 5'h17 == csrs_8_Index ? tlb_23_P1_PLV : _GEN_664;
  wire [1:0] _GEN_666 = 5'h18 == csrs_8_Index ? tlb_24_P1_PLV : _GEN_665;
  wire [1:0] _GEN_667 = 5'h19 == csrs_8_Index ? tlb_25_P1_PLV : _GEN_666;
  wire [1:0] _GEN_668 = 5'h1a == csrs_8_Index ? tlb_26_P1_PLV : _GEN_667;
  wire [1:0] _GEN_669 = 5'h1b == csrs_8_Index ? tlb_27_P1_PLV : _GEN_668;
  wire [1:0] _GEN_670 = 5'h1c == csrs_8_Index ? tlb_28_P1_PLV : _GEN_669;
  wire [1:0] _GEN_671 = 5'h1d == csrs_8_Index ? tlb_29_P1_PLV : _GEN_670;
  wire [1:0] _GEN_672 = 5'h1e == csrs_8_Index ? tlb_30_P1_PLV : _GEN_671;
  wire [1:0] _GEN_673 = 5'h1f == csrs_8_Index ? tlb_31_P1_PLV : _GEN_672;
  wire  _GEN_675 = 5'h1 == csrs_8_Index ? tlb_1_P1_D : tlb_0_P1_D;
  wire  _GEN_676 = 5'h2 == csrs_8_Index ? tlb_2_P1_D : _GEN_675;
  wire  _GEN_677 = 5'h3 == csrs_8_Index ? tlb_3_P1_D : _GEN_676;
  wire  _GEN_678 = 5'h4 == csrs_8_Index ? tlb_4_P1_D : _GEN_677;
  wire  _GEN_679 = 5'h5 == csrs_8_Index ? tlb_5_P1_D : _GEN_678;
  wire  _GEN_680 = 5'h6 == csrs_8_Index ? tlb_6_P1_D : _GEN_679;
  wire  _GEN_681 = 5'h7 == csrs_8_Index ? tlb_7_P1_D : _GEN_680;
  wire  _GEN_682 = 5'h8 == csrs_8_Index ? tlb_8_P1_D : _GEN_681;
  wire  _GEN_683 = 5'h9 == csrs_8_Index ? tlb_9_P1_D : _GEN_682;
  wire  _GEN_684 = 5'ha == csrs_8_Index ? tlb_10_P1_D : _GEN_683;
  wire  _GEN_685 = 5'hb == csrs_8_Index ? tlb_11_P1_D : _GEN_684;
  wire  _GEN_686 = 5'hc == csrs_8_Index ? tlb_12_P1_D : _GEN_685;
  wire  _GEN_687 = 5'hd == csrs_8_Index ? tlb_13_P1_D : _GEN_686;
  wire  _GEN_688 = 5'he == csrs_8_Index ? tlb_14_P1_D : _GEN_687;
  wire  _GEN_689 = 5'hf == csrs_8_Index ? tlb_15_P1_D : _GEN_688;
  wire  _GEN_690 = 5'h10 == csrs_8_Index ? tlb_16_P1_D : _GEN_689;
  wire  _GEN_691 = 5'h11 == csrs_8_Index ? tlb_17_P1_D : _GEN_690;
  wire  _GEN_692 = 5'h12 == csrs_8_Index ? tlb_18_P1_D : _GEN_691;
  wire  _GEN_693 = 5'h13 == csrs_8_Index ? tlb_19_P1_D : _GEN_692;
  wire  _GEN_694 = 5'h14 == csrs_8_Index ? tlb_20_P1_D : _GEN_693;
  wire  _GEN_695 = 5'h15 == csrs_8_Index ? tlb_21_P1_D : _GEN_694;
  wire  _GEN_696 = 5'h16 == csrs_8_Index ? tlb_22_P1_D : _GEN_695;
  wire  _GEN_697 = 5'h17 == csrs_8_Index ? tlb_23_P1_D : _GEN_696;
  wire  _GEN_698 = 5'h18 == csrs_8_Index ? tlb_24_P1_D : _GEN_697;
  wire  _GEN_699 = 5'h19 == csrs_8_Index ? tlb_25_P1_D : _GEN_698;
  wire  _GEN_700 = 5'h1a == csrs_8_Index ? tlb_26_P1_D : _GEN_699;
  wire  _GEN_701 = 5'h1b == csrs_8_Index ? tlb_27_P1_D : _GEN_700;
  wire  _GEN_702 = 5'h1c == csrs_8_Index ? tlb_28_P1_D : _GEN_701;
  wire  _GEN_703 = 5'h1d == csrs_8_Index ? tlb_29_P1_D : _GEN_702;
  wire  _GEN_704 = 5'h1e == csrs_8_Index ? tlb_30_P1_D : _GEN_703;
  wire  _GEN_705 = 5'h1f == csrs_8_Index ? tlb_31_P1_D : _GEN_704;
  wire  _GEN_707 = 5'h1 == csrs_8_Index ? tlb_1_P1_V : tlb_0_P1_V;
  wire  _GEN_708 = 5'h2 == csrs_8_Index ? tlb_2_P1_V : _GEN_707;
  wire  _GEN_709 = 5'h3 == csrs_8_Index ? tlb_3_P1_V : _GEN_708;
  wire  _GEN_710 = 5'h4 == csrs_8_Index ? tlb_4_P1_V : _GEN_709;
  wire  _GEN_711 = 5'h5 == csrs_8_Index ? tlb_5_P1_V : _GEN_710;
  wire  _GEN_712 = 5'h6 == csrs_8_Index ? tlb_6_P1_V : _GEN_711;
  wire  _GEN_713 = 5'h7 == csrs_8_Index ? tlb_7_P1_V : _GEN_712;
  wire  _GEN_714 = 5'h8 == csrs_8_Index ? tlb_8_P1_V : _GEN_713;
  wire  _GEN_715 = 5'h9 == csrs_8_Index ? tlb_9_P1_V : _GEN_714;
  wire  _GEN_716 = 5'ha == csrs_8_Index ? tlb_10_P1_V : _GEN_715;
  wire  _GEN_717 = 5'hb == csrs_8_Index ? tlb_11_P1_V : _GEN_716;
  wire  _GEN_718 = 5'hc == csrs_8_Index ? tlb_12_P1_V : _GEN_717;
  wire  _GEN_719 = 5'hd == csrs_8_Index ? tlb_13_P1_V : _GEN_718;
  wire  _GEN_720 = 5'he == csrs_8_Index ? tlb_14_P1_V : _GEN_719;
  wire  _GEN_721 = 5'hf == csrs_8_Index ? tlb_15_P1_V : _GEN_720;
  wire  _GEN_722 = 5'h10 == csrs_8_Index ? tlb_16_P1_V : _GEN_721;
  wire  _GEN_723 = 5'h11 == csrs_8_Index ? tlb_17_P1_V : _GEN_722;
  wire  _GEN_724 = 5'h12 == csrs_8_Index ? tlb_18_P1_V : _GEN_723;
  wire  _GEN_725 = 5'h13 == csrs_8_Index ? tlb_19_P1_V : _GEN_724;
  wire  _GEN_726 = 5'h14 == csrs_8_Index ? tlb_20_P1_V : _GEN_725;
  wire  _GEN_727 = 5'h15 == csrs_8_Index ? tlb_21_P1_V : _GEN_726;
  wire  _GEN_728 = 5'h16 == csrs_8_Index ? tlb_22_P1_V : _GEN_727;
  wire  _GEN_729 = 5'h17 == csrs_8_Index ? tlb_23_P1_V : _GEN_728;
  wire  _GEN_730 = 5'h18 == csrs_8_Index ? tlb_24_P1_V : _GEN_729;
  wire  _GEN_731 = 5'h19 == csrs_8_Index ? tlb_25_P1_V : _GEN_730;
  wire  _GEN_732 = 5'h1a == csrs_8_Index ? tlb_26_P1_V : _GEN_731;
  wire  _GEN_733 = 5'h1b == csrs_8_Index ? tlb_27_P1_V : _GEN_732;
  wire  _GEN_734 = 5'h1c == csrs_8_Index ? tlb_28_P1_V : _GEN_733;
  wire  _GEN_735 = 5'h1d == csrs_8_Index ? tlb_29_P1_V : _GEN_734;
  wire  _GEN_736 = 5'h1e == csrs_8_Index ? tlb_30_P1_V : _GEN_735;
  wire  _GEN_737 = 5'h1f == csrs_8_Index ? tlb_31_P1_V : _GEN_736;
  wire [9:0] _GEN_739 = 5'h1 == csrs_8_Index ? tlb_1_ASID : tlb_0_ASID;
  wire [9:0] _GEN_740 = 5'h2 == csrs_8_Index ? tlb_2_ASID : _GEN_739;
  wire [9:0] _GEN_741 = 5'h3 == csrs_8_Index ? tlb_3_ASID : _GEN_740;
  wire [9:0] _GEN_742 = 5'h4 == csrs_8_Index ? tlb_4_ASID : _GEN_741;
  wire [9:0] _GEN_743 = 5'h5 == csrs_8_Index ? tlb_5_ASID : _GEN_742;
  wire [9:0] _GEN_744 = 5'h6 == csrs_8_Index ? tlb_6_ASID : _GEN_743;
  wire [9:0] _GEN_745 = 5'h7 == csrs_8_Index ? tlb_7_ASID : _GEN_744;
  wire [9:0] _GEN_746 = 5'h8 == csrs_8_Index ? tlb_8_ASID : _GEN_745;
  wire [9:0] _GEN_747 = 5'h9 == csrs_8_Index ? tlb_9_ASID : _GEN_746;
  wire [9:0] _GEN_748 = 5'ha == csrs_8_Index ? tlb_10_ASID : _GEN_747;
  wire [9:0] _GEN_749 = 5'hb == csrs_8_Index ? tlb_11_ASID : _GEN_748;
  wire [9:0] _GEN_750 = 5'hc == csrs_8_Index ? tlb_12_ASID : _GEN_749;
  wire [9:0] _GEN_751 = 5'hd == csrs_8_Index ? tlb_13_ASID : _GEN_750;
  wire [9:0] _GEN_752 = 5'he == csrs_8_Index ? tlb_14_ASID : _GEN_751;
  wire [9:0] _GEN_753 = 5'hf == csrs_8_Index ? tlb_15_ASID : _GEN_752;
  wire [9:0] _GEN_754 = 5'h10 == csrs_8_Index ? tlb_16_ASID : _GEN_753;
  wire [9:0] _GEN_755 = 5'h11 == csrs_8_Index ? tlb_17_ASID : _GEN_754;
  wire [9:0] _GEN_756 = 5'h12 == csrs_8_Index ? tlb_18_ASID : _GEN_755;
  wire [9:0] _GEN_757 = 5'h13 == csrs_8_Index ? tlb_19_ASID : _GEN_756;
  wire [9:0] _GEN_758 = 5'h14 == csrs_8_Index ? tlb_20_ASID : _GEN_757;
  wire [9:0] _GEN_759 = 5'h15 == csrs_8_Index ? tlb_21_ASID : _GEN_758;
  wire [9:0] _GEN_760 = 5'h16 == csrs_8_Index ? tlb_22_ASID : _GEN_759;
  wire [9:0] _GEN_761 = 5'h17 == csrs_8_Index ? tlb_23_ASID : _GEN_760;
  wire [9:0] _GEN_762 = 5'h18 == csrs_8_Index ? tlb_24_ASID : _GEN_761;
  wire [9:0] _GEN_763 = 5'h19 == csrs_8_Index ? tlb_25_ASID : _GEN_762;
  wire [9:0] _GEN_764 = 5'h1a == csrs_8_Index ? tlb_26_ASID : _GEN_763;
  wire [9:0] _GEN_765 = 5'h1b == csrs_8_Index ? tlb_27_ASID : _GEN_764;
  wire [9:0] _GEN_766 = 5'h1c == csrs_8_Index ? tlb_28_ASID : _GEN_765;
  wire [9:0] _GEN_767 = 5'h1d == csrs_8_Index ? tlb_29_ASID : _GEN_766;
  wire [9:0] _GEN_768 = 5'h1e == csrs_8_Index ? tlb_30_ASID : _GEN_767;
  wire [9:0] _GEN_769 = 5'h1f == csrs_8_Index ? tlb_31_ASID : _GEN_768;
  wire [5:0] _GEN_770 = _GEN_321 ? _GEN_353 : _GEN_247;
  wire [18:0] _GEN_771 = _GEN_321 ? _GEN_385 : _GEN_249;
  wire [23:0] _GEN_772 = _GEN_321 ? {{4'd0}, _GEN_417} : _GEN_255;
  wire  _GEN_773 = _GEN_321 ? _GEN_449 : _GEN_254;
  wire [1:0] _GEN_774 = _GEN_321 ? _GEN_481 : _GEN_253;
  wire [1:0] _GEN_775 = _GEN_321 ? _GEN_513 : _GEN_252;
  wire  _GEN_776 = _GEN_321 ? _GEN_545 : _GEN_251;
  wire  _GEN_777 = _GEN_321 ? _GEN_577 : _GEN_250;
  wire [23:0] _GEN_778 = _GEN_321 ? {{4'd0}, _GEN_609} : _GEN_261;
  wire  _GEN_779 = _GEN_321 ? _GEN_449 : _GEN_260;
  wire [1:0] _GEN_780 = _GEN_321 ? _GEN_641 : _GEN_259;
  wire [1:0] _GEN_781 = _GEN_321 ? _GEN_673 : _GEN_258;
  wire  _GEN_782 = _GEN_321 ? _GEN_705 : _GEN_257;
  wire  _GEN_783 = _GEN_321 ? _GEN_737 : _GEN_256;
  wire [9:0] _GEN_784 = _GEN_321 ? _GEN_769 : _GEN_262;
  wire [18:0] _GEN_785 = 5'h0 == csrs_8_Index ? csrs_9_VPPN : tlb_0_VPPN;
  wire [18:0] _GEN_786 = 5'h1 == csrs_8_Index ? csrs_9_VPPN : tlb_1_VPPN;
  wire [18:0] _GEN_787 = 5'h2 == csrs_8_Index ? csrs_9_VPPN : tlb_2_VPPN;
  wire [18:0] _GEN_788 = 5'h3 == csrs_8_Index ? csrs_9_VPPN : tlb_3_VPPN;
  wire [18:0] _GEN_789 = 5'h4 == csrs_8_Index ? csrs_9_VPPN : tlb_4_VPPN;
  wire [18:0] _GEN_790 = 5'h5 == csrs_8_Index ? csrs_9_VPPN : tlb_5_VPPN;
  wire [18:0] _GEN_791 = 5'h6 == csrs_8_Index ? csrs_9_VPPN : tlb_6_VPPN;
  wire [18:0] _GEN_792 = 5'h7 == csrs_8_Index ? csrs_9_VPPN : tlb_7_VPPN;
  wire [18:0] _GEN_793 = 5'h8 == csrs_8_Index ? csrs_9_VPPN : tlb_8_VPPN;
  wire [18:0] _GEN_794 = 5'h9 == csrs_8_Index ? csrs_9_VPPN : tlb_9_VPPN;
  wire [18:0] _GEN_795 = 5'ha == csrs_8_Index ? csrs_9_VPPN : tlb_10_VPPN;
  wire [18:0] _GEN_796 = 5'hb == csrs_8_Index ? csrs_9_VPPN : tlb_11_VPPN;
  wire [18:0] _GEN_797 = 5'hc == csrs_8_Index ? csrs_9_VPPN : tlb_12_VPPN;
  wire [18:0] _GEN_798 = 5'hd == csrs_8_Index ? csrs_9_VPPN : tlb_13_VPPN;
  wire [18:0] _GEN_799 = 5'he == csrs_8_Index ? csrs_9_VPPN : tlb_14_VPPN;
  wire [18:0] _GEN_800 = 5'hf == csrs_8_Index ? csrs_9_VPPN : tlb_15_VPPN;
  wire [18:0] _GEN_801 = 5'h10 == csrs_8_Index ? csrs_9_VPPN : tlb_16_VPPN;
  wire [18:0] _GEN_802 = 5'h11 == csrs_8_Index ? csrs_9_VPPN : tlb_17_VPPN;
  wire [18:0] _GEN_803 = 5'h12 == csrs_8_Index ? csrs_9_VPPN : tlb_18_VPPN;
  wire [18:0] _GEN_804 = 5'h13 == csrs_8_Index ? csrs_9_VPPN : tlb_19_VPPN;
  wire [18:0] _GEN_805 = 5'h14 == csrs_8_Index ? csrs_9_VPPN : tlb_20_VPPN;
  wire [18:0] _GEN_806 = 5'h15 == csrs_8_Index ? csrs_9_VPPN : tlb_21_VPPN;
  wire [18:0] _GEN_807 = 5'h16 == csrs_8_Index ? csrs_9_VPPN : tlb_22_VPPN;
  wire [18:0] _GEN_808 = 5'h17 == csrs_8_Index ? csrs_9_VPPN : tlb_23_VPPN;
  wire [18:0] _GEN_809 = 5'h18 == csrs_8_Index ? csrs_9_VPPN : tlb_24_VPPN;
  wire [18:0] _GEN_810 = 5'h19 == csrs_8_Index ? csrs_9_VPPN : tlb_25_VPPN;
  wire [18:0] _GEN_811 = 5'h1a == csrs_8_Index ? csrs_9_VPPN : tlb_26_VPPN;
  wire [18:0] _GEN_812 = 5'h1b == csrs_8_Index ? csrs_9_VPPN : tlb_27_VPPN;
  wire [18:0] _GEN_813 = 5'h1c == csrs_8_Index ? csrs_9_VPPN : tlb_28_VPPN;
  wire [18:0] _GEN_814 = 5'h1d == csrs_8_Index ? csrs_9_VPPN : tlb_29_VPPN;
  wire [18:0] _GEN_815 = 5'h1e == csrs_8_Index ? csrs_9_VPPN : tlb_30_VPPN;
  wire [18:0] _GEN_816 = 5'h1f == csrs_8_Index ? csrs_9_VPPN : tlb_31_VPPN;
  wire [5:0] _GEN_817 = 5'h0 == csrs_8_Index ? csrs_8_PS : tlb_0_PS;
  wire [5:0] _GEN_818 = 5'h1 == csrs_8_Index ? csrs_8_PS : tlb_1_PS;
  wire [5:0] _GEN_819 = 5'h2 == csrs_8_Index ? csrs_8_PS : tlb_2_PS;
  wire [5:0] _GEN_820 = 5'h3 == csrs_8_Index ? csrs_8_PS : tlb_3_PS;
  wire [5:0] _GEN_821 = 5'h4 == csrs_8_Index ? csrs_8_PS : tlb_4_PS;
  wire [5:0] _GEN_822 = 5'h5 == csrs_8_Index ? csrs_8_PS : tlb_5_PS;
  wire [5:0] _GEN_823 = 5'h6 == csrs_8_Index ? csrs_8_PS : tlb_6_PS;
  wire [5:0] _GEN_824 = 5'h7 == csrs_8_Index ? csrs_8_PS : tlb_7_PS;
  wire [5:0] _GEN_825 = 5'h8 == csrs_8_Index ? csrs_8_PS : tlb_8_PS;
  wire [5:0] _GEN_826 = 5'h9 == csrs_8_Index ? csrs_8_PS : tlb_9_PS;
  wire [5:0] _GEN_827 = 5'ha == csrs_8_Index ? csrs_8_PS : tlb_10_PS;
  wire [5:0] _GEN_828 = 5'hb == csrs_8_Index ? csrs_8_PS : tlb_11_PS;
  wire [5:0] _GEN_829 = 5'hc == csrs_8_Index ? csrs_8_PS : tlb_12_PS;
  wire [5:0] _GEN_830 = 5'hd == csrs_8_Index ? csrs_8_PS : tlb_13_PS;
  wire [5:0] _GEN_831 = 5'he == csrs_8_Index ? csrs_8_PS : tlb_14_PS;
  wire [5:0] _GEN_832 = 5'hf == csrs_8_Index ? csrs_8_PS : tlb_15_PS;
  wire [5:0] _GEN_833 = 5'h10 == csrs_8_Index ? csrs_8_PS : tlb_16_PS;
  wire [5:0] _GEN_834 = 5'h11 == csrs_8_Index ? csrs_8_PS : tlb_17_PS;
  wire [5:0] _GEN_835 = 5'h12 == csrs_8_Index ? csrs_8_PS : tlb_18_PS;
  wire [5:0] _GEN_836 = 5'h13 == csrs_8_Index ? csrs_8_PS : tlb_19_PS;
  wire [5:0] _GEN_837 = 5'h14 == csrs_8_Index ? csrs_8_PS : tlb_20_PS;
  wire [5:0] _GEN_838 = 5'h15 == csrs_8_Index ? csrs_8_PS : tlb_21_PS;
  wire [5:0] _GEN_839 = 5'h16 == csrs_8_Index ? csrs_8_PS : tlb_22_PS;
  wire [5:0] _GEN_840 = 5'h17 == csrs_8_Index ? csrs_8_PS : tlb_23_PS;
  wire [5:0] _GEN_841 = 5'h18 == csrs_8_Index ? csrs_8_PS : tlb_24_PS;
  wire [5:0] _GEN_842 = 5'h19 == csrs_8_Index ? csrs_8_PS : tlb_25_PS;
  wire [5:0] _GEN_843 = 5'h1a == csrs_8_Index ? csrs_8_PS : tlb_26_PS;
  wire [5:0] _GEN_844 = 5'h1b == csrs_8_Index ? csrs_8_PS : tlb_27_PS;
  wire [5:0] _GEN_845 = 5'h1c == csrs_8_Index ? csrs_8_PS : tlb_28_PS;
  wire [5:0] _GEN_846 = 5'h1d == csrs_8_Index ? csrs_8_PS : tlb_29_PS;
  wire [5:0] _GEN_847 = 5'h1e == csrs_8_Index ? csrs_8_PS : tlb_30_PS;
  wire [5:0] _GEN_848 = 5'h1f == csrs_8_Index ? csrs_8_PS : tlb_31_PS;
  wire  _GEN_849 = 5'h0 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_0_G;
  wire  _GEN_850 = 5'h1 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_1_G;
  wire  _GEN_851 = 5'h2 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_2_G;
  wire  _GEN_852 = 5'h3 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_3_G;
  wire  _GEN_853 = 5'h4 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_4_G;
  wire  _GEN_854 = 5'h5 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_5_G;
  wire  _GEN_855 = 5'h6 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_6_G;
  wire  _GEN_856 = 5'h7 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_7_G;
  wire  _GEN_857 = 5'h8 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_8_G;
  wire  _GEN_858 = 5'h9 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_9_G;
  wire  _GEN_859 = 5'ha == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_10_G;
  wire  _GEN_860 = 5'hb == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_11_G;
  wire  _GEN_861 = 5'hc == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_12_G;
  wire  _GEN_862 = 5'hd == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_13_G;
  wire  _GEN_863 = 5'he == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_14_G;
  wire  _GEN_864 = 5'hf == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_15_G;
  wire  _GEN_865 = 5'h10 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_16_G;
  wire  _GEN_866 = 5'h11 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_17_G;
  wire  _GEN_867 = 5'h12 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_18_G;
  wire  _GEN_868 = 5'h13 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_19_G;
  wire  _GEN_869 = 5'h14 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_20_G;
  wire  _GEN_870 = 5'h15 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_21_G;
  wire  _GEN_871 = 5'h16 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_22_G;
  wire  _GEN_872 = 5'h17 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_23_G;
  wire  _GEN_873 = 5'h18 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_24_G;
  wire  _GEN_874 = 5'h19 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_25_G;
  wire  _GEN_875 = 5'h1a == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_26_G;
  wire  _GEN_876 = 5'h1b == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_27_G;
  wire  _GEN_877 = 5'h1c == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_28_G;
  wire  _GEN_878 = 5'h1d == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_29_G;
  wire  _GEN_879 = 5'h1e == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_30_G;
  wire  _GEN_880 = 5'h1f == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_31_G;
  wire [9:0] _GEN_881 = 5'h0 == csrs_8_Index ? asid_ASID : tlb_0_ASID;
  wire [9:0] _GEN_882 = 5'h1 == csrs_8_Index ? asid_ASID : tlb_1_ASID;
  wire [9:0] _GEN_883 = 5'h2 == csrs_8_Index ? asid_ASID : tlb_2_ASID;
  wire [9:0] _GEN_884 = 5'h3 == csrs_8_Index ? asid_ASID : tlb_3_ASID;
  wire [9:0] _GEN_885 = 5'h4 == csrs_8_Index ? asid_ASID : tlb_4_ASID;
  wire [9:0] _GEN_886 = 5'h5 == csrs_8_Index ? asid_ASID : tlb_5_ASID;
  wire [9:0] _GEN_887 = 5'h6 == csrs_8_Index ? asid_ASID : tlb_6_ASID;
  wire [9:0] _GEN_888 = 5'h7 == csrs_8_Index ? asid_ASID : tlb_7_ASID;
  wire [9:0] _GEN_889 = 5'h8 == csrs_8_Index ? asid_ASID : tlb_8_ASID;
  wire [9:0] _GEN_890 = 5'h9 == csrs_8_Index ? asid_ASID : tlb_9_ASID;
  wire [9:0] _GEN_891 = 5'ha == csrs_8_Index ? asid_ASID : tlb_10_ASID;
  wire [9:0] _GEN_892 = 5'hb == csrs_8_Index ? asid_ASID : tlb_11_ASID;
  wire [9:0] _GEN_893 = 5'hc == csrs_8_Index ? asid_ASID : tlb_12_ASID;
  wire [9:0] _GEN_894 = 5'hd == csrs_8_Index ? asid_ASID : tlb_13_ASID;
  wire [9:0] _GEN_895 = 5'he == csrs_8_Index ? asid_ASID : tlb_14_ASID;
  wire [9:0] _GEN_896 = 5'hf == csrs_8_Index ? asid_ASID : tlb_15_ASID;
  wire [9:0] _GEN_897 = 5'h10 == csrs_8_Index ? asid_ASID : tlb_16_ASID;
  wire [9:0] _GEN_898 = 5'h11 == csrs_8_Index ? asid_ASID : tlb_17_ASID;
  wire [9:0] _GEN_899 = 5'h12 == csrs_8_Index ? asid_ASID : tlb_18_ASID;
  wire [9:0] _GEN_900 = 5'h13 == csrs_8_Index ? asid_ASID : tlb_19_ASID;
  wire [9:0] _GEN_901 = 5'h14 == csrs_8_Index ? asid_ASID : tlb_20_ASID;
  wire [9:0] _GEN_902 = 5'h15 == csrs_8_Index ? asid_ASID : tlb_21_ASID;
  wire [9:0] _GEN_903 = 5'h16 == csrs_8_Index ? asid_ASID : tlb_22_ASID;
  wire [9:0] _GEN_904 = 5'h17 == csrs_8_Index ? asid_ASID : tlb_23_ASID;
  wire [9:0] _GEN_905 = 5'h18 == csrs_8_Index ? asid_ASID : tlb_24_ASID;
  wire [9:0] _GEN_906 = 5'h19 == csrs_8_Index ? asid_ASID : tlb_25_ASID;
  wire [9:0] _GEN_907 = 5'h1a == csrs_8_Index ? asid_ASID : tlb_26_ASID;
  wire [9:0] _GEN_908 = 5'h1b == csrs_8_Index ? asid_ASID : tlb_27_ASID;
  wire [9:0] _GEN_909 = 5'h1c == csrs_8_Index ? asid_ASID : tlb_28_ASID;
  wire [9:0] _GEN_910 = 5'h1d == csrs_8_Index ? asid_ASID : tlb_29_ASID;
  wire [9:0] _GEN_911 = 5'h1e == csrs_8_Index ? asid_ASID : tlb_30_ASID;
  wire [9:0] _GEN_912 = 5'h1f == csrs_8_Index ? asid_ASID : tlb_31_ASID;
  wire  _tlb_E_T = csrs_4_Ecode == 6'h3f;
  wire  _GEN_913 = 5'h0 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_0_E;
  wire  _GEN_914 = 5'h1 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_1_E;
  wire  _GEN_915 = 5'h2 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_2_E;
  wire  _GEN_916 = 5'h3 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_3_E;
  wire  _GEN_917 = 5'h4 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_4_E;
  wire  _GEN_918 = 5'h5 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_5_E;
  wire  _GEN_919 = 5'h6 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_6_E;
  wire  _GEN_920 = 5'h7 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_7_E;
  wire  _GEN_921 = 5'h8 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_8_E;
  wire  _GEN_922 = 5'h9 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_9_E;
  wire  _GEN_923 = 5'ha == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_10_E;
  wire  _GEN_924 = 5'hb == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_11_E;
  wire  _GEN_925 = 5'hc == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_12_E;
  wire  _GEN_926 = 5'hd == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_13_E;
  wire  _GEN_927 = 5'he == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_14_E;
  wire  _GEN_928 = 5'hf == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_15_E;
  wire  _GEN_929 = 5'h10 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_16_E;
  wire  _GEN_930 = 5'h11 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_17_E;
  wire  _GEN_931 = 5'h12 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_18_E;
  wire  _GEN_932 = 5'h13 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_19_E;
  wire  _GEN_933 = 5'h14 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_20_E;
  wire  _GEN_934 = 5'h15 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_21_E;
  wire  _GEN_935 = 5'h16 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_22_E;
  wire  _GEN_936 = 5'h17 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_23_E;
  wire  _GEN_937 = 5'h18 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_24_E;
  wire  _GEN_938 = 5'h19 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_25_E;
  wire  _GEN_939 = 5'h1a == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_26_E;
  wire  _GEN_940 = 5'h1b == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_27_E;
  wire  _GEN_941 = 5'h1c == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_28_E;
  wire  _GEN_942 = 5'h1d == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_29_E;
  wire  _GEN_943 = 5'h1e == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_30_E;
  wire  _GEN_944 = 5'h1f == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_31_E;
  wire [19:0] _GEN_945 = 5'h0 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_0_P0_PPN;
  wire [19:0] _GEN_946 = 5'h1 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_1_P0_PPN;
  wire [19:0] _GEN_947 = 5'h2 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_2_P0_PPN;
  wire [19:0] _GEN_948 = 5'h3 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_3_P0_PPN;
  wire [19:0] _GEN_949 = 5'h4 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_4_P0_PPN;
  wire [19:0] _GEN_950 = 5'h5 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_5_P0_PPN;
  wire [19:0] _GEN_951 = 5'h6 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_6_P0_PPN;
  wire [19:0] _GEN_952 = 5'h7 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_7_P0_PPN;
  wire [19:0] _GEN_953 = 5'h8 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_8_P0_PPN;
  wire [19:0] _GEN_954 = 5'h9 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_9_P0_PPN;
  wire [19:0] _GEN_955 = 5'ha == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_10_P0_PPN;
  wire [19:0] _GEN_956 = 5'hb == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_11_P0_PPN;
  wire [19:0] _GEN_957 = 5'hc == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_12_P0_PPN;
  wire [19:0] _GEN_958 = 5'hd == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_13_P0_PPN;
  wire [19:0] _GEN_959 = 5'he == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_14_P0_PPN;
  wire [19:0] _GEN_960 = 5'hf == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_15_P0_PPN;
  wire [19:0] _GEN_961 = 5'h10 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_16_P0_PPN;
  wire [19:0] _GEN_962 = 5'h11 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_17_P0_PPN;
  wire [19:0] _GEN_963 = 5'h12 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_18_P0_PPN;
  wire [19:0] _GEN_964 = 5'h13 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_19_P0_PPN;
  wire [19:0] _GEN_965 = 5'h14 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_20_P0_PPN;
  wire [19:0] _GEN_966 = 5'h15 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_21_P0_PPN;
  wire [19:0] _GEN_967 = 5'h16 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_22_P0_PPN;
  wire [19:0] _GEN_968 = 5'h17 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_23_P0_PPN;
  wire [19:0] _GEN_969 = 5'h18 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_24_P0_PPN;
  wire [19:0] _GEN_970 = 5'h19 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_25_P0_PPN;
  wire [19:0] _GEN_971 = 5'h1a == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_26_P0_PPN;
  wire [19:0] _GEN_972 = 5'h1b == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_27_P0_PPN;
  wire [19:0] _GEN_973 = 5'h1c == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_28_P0_PPN;
  wire [19:0] _GEN_974 = 5'h1d == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_29_P0_PPN;
  wire [19:0] _GEN_975 = 5'h1e == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_30_P0_PPN;
  wire [19:0] _GEN_976 = 5'h1f == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_31_P0_PPN;
  wire [1:0] _GEN_977 = 5'h0 == csrs_8_Index ? csrs_10_PLV : tlb_0_P0_PLV;
  wire [1:0] _GEN_978 = 5'h1 == csrs_8_Index ? csrs_10_PLV : tlb_1_P0_PLV;
  wire [1:0] _GEN_979 = 5'h2 == csrs_8_Index ? csrs_10_PLV : tlb_2_P0_PLV;
  wire [1:0] _GEN_980 = 5'h3 == csrs_8_Index ? csrs_10_PLV : tlb_3_P0_PLV;
  wire [1:0] _GEN_981 = 5'h4 == csrs_8_Index ? csrs_10_PLV : tlb_4_P0_PLV;
  wire [1:0] _GEN_982 = 5'h5 == csrs_8_Index ? csrs_10_PLV : tlb_5_P0_PLV;
  wire [1:0] _GEN_983 = 5'h6 == csrs_8_Index ? csrs_10_PLV : tlb_6_P0_PLV;
  wire [1:0] _GEN_984 = 5'h7 == csrs_8_Index ? csrs_10_PLV : tlb_7_P0_PLV;
  wire [1:0] _GEN_985 = 5'h8 == csrs_8_Index ? csrs_10_PLV : tlb_8_P0_PLV;
  wire [1:0] _GEN_986 = 5'h9 == csrs_8_Index ? csrs_10_PLV : tlb_9_P0_PLV;
  wire [1:0] _GEN_987 = 5'ha == csrs_8_Index ? csrs_10_PLV : tlb_10_P0_PLV;
  wire [1:0] _GEN_988 = 5'hb == csrs_8_Index ? csrs_10_PLV : tlb_11_P0_PLV;
  wire [1:0] _GEN_989 = 5'hc == csrs_8_Index ? csrs_10_PLV : tlb_12_P0_PLV;
  wire [1:0] _GEN_990 = 5'hd == csrs_8_Index ? csrs_10_PLV : tlb_13_P0_PLV;
  wire [1:0] _GEN_991 = 5'he == csrs_8_Index ? csrs_10_PLV : tlb_14_P0_PLV;
  wire [1:0] _GEN_992 = 5'hf == csrs_8_Index ? csrs_10_PLV : tlb_15_P0_PLV;
  wire [1:0] _GEN_993 = 5'h10 == csrs_8_Index ? csrs_10_PLV : tlb_16_P0_PLV;
  wire [1:0] _GEN_994 = 5'h11 == csrs_8_Index ? csrs_10_PLV : tlb_17_P0_PLV;
  wire [1:0] _GEN_995 = 5'h12 == csrs_8_Index ? csrs_10_PLV : tlb_18_P0_PLV;
  wire [1:0] _GEN_996 = 5'h13 == csrs_8_Index ? csrs_10_PLV : tlb_19_P0_PLV;
  wire [1:0] _GEN_997 = 5'h14 == csrs_8_Index ? csrs_10_PLV : tlb_20_P0_PLV;
  wire [1:0] _GEN_998 = 5'h15 == csrs_8_Index ? csrs_10_PLV : tlb_21_P0_PLV;
  wire [1:0] _GEN_999 = 5'h16 == csrs_8_Index ? csrs_10_PLV : tlb_22_P0_PLV;
  wire [1:0] _GEN_1000 = 5'h17 == csrs_8_Index ? csrs_10_PLV : tlb_23_P0_PLV;
  wire [1:0] _GEN_1001 = 5'h18 == csrs_8_Index ? csrs_10_PLV : tlb_24_P0_PLV;
  wire [1:0] _GEN_1002 = 5'h19 == csrs_8_Index ? csrs_10_PLV : tlb_25_P0_PLV;
  wire [1:0] _GEN_1003 = 5'h1a == csrs_8_Index ? csrs_10_PLV : tlb_26_P0_PLV;
  wire [1:0] _GEN_1004 = 5'h1b == csrs_8_Index ? csrs_10_PLV : tlb_27_P0_PLV;
  wire [1:0] _GEN_1005 = 5'h1c == csrs_8_Index ? csrs_10_PLV : tlb_28_P0_PLV;
  wire [1:0] _GEN_1006 = 5'h1d == csrs_8_Index ? csrs_10_PLV : tlb_29_P0_PLV;
  wire [1:0] _GEN_1007 = 5'h1e == csrs_8_Index ? csrs_10_PLV : tlb_30_P0_PLV;
  wire [1:0] _GEN_1008 = 5'h1f == csrs_8_Index ? csrs_10_PLV : tlb_31_P0_PLV;
  wire [1:0] _GEN_1009 = 5'h0 == csrs_8_Index ? csrs_10_MAT : tlb_0_P0_MAT;
  wire [1:0] _GEN_1010 = 5'h1 == csrs_8_Index ? csrs_10_MAT : tlb_1_P0_MAT;
  wire [1:0] _GEN_1011 = 5'h2 == csrs_8_Index ? csrs_10_MAT : tlb_2_P0_MAT;
  wire [1:0] _GEN_1012 = 5'h3 == csrs_8_Index ? csrs_10_MAT : tlb_3_P0_MAT;
  wire [1:0] _GEN_1013 = 5'h4 == csrs_8_Index ? csrs_10_MAT : tlb_4_P0_MAT;
  wire [1:0] _GEN_1014 = 5'h5 == csrs_8_Index ? csrs_10_MAT : tlb_5_P0_MAT;
  wire [1:0] _GEN_1015 = 5'h6 == csrs_8_Index ? csrs_10_MAT : tlb_6_P0_MAT;
  wire [1:0] _GEN_1016 = 5'h7 == csrs_8_Index ? csrs_10_MAT : tlb_7_P0_MAT;
  wire [1:0] _GEN_1017 = 5'h8 == csrs_8_Index ? csrs_10_MAT : tlb_8_P0_MAT;
  wire [1:0] _GEN_1018 = 5'h9 == csrs_8_Index ? csrs_10_MAT : tlb_9_P0_MAT;
  wire [1:0] _GEN_1019 = 5'ha == csrs_8_Index ? csrs_10_MAT : tlb_10_P0_MAT;
  wire [1:0] _GEN_1020 = 5'hb == csrs_8_Index ? csrs_10_MAT : tlb_11_P0_MAT;
  wire [1:0] _GEN_1021 = 5'hc == csrs_8_Index ? csrs_10_MAT : tlb_12_P0_MAT;
  wire [1:0] _GEN_1022 = 5'hd == csrs_8_Index ? csrs_10_MAT : tlb_13_P0_MAT;
  wire [1:0] _GEN_1023 = 5'he == csrs_8_Index ? csrs_10_MAT : tlb_14_P0_MAT;
  wire [1:0] _GEN_1024 = 5'hf == csrs_8_Index ? csrs_10_MAT : tlb_15_P0_MAT;
  wire [1:0] _GEN_1025 = 5'h10 == csrs_8_Index ? csrs_10_MAT : tlb_16_P0_MAT;
  wire [1:0] _GEN_1026 = 5'h11 == csrs_8_Index ? csrs_10_MAT : tlb_17_P0_MAT;
  wire [1:0] _GEN_1027 = 5'h12 == csrs_8_Index ? csrs_10_MAT : tlb_18_P0_MAT;
  wire [1:0] _GEN_1028 = 5'h13 == csrs_8_Index ? csrs_10_MAT : tlb_19_P0_MAT;
  wire [1:0] _GEN_1029 = 5'h14 == csrs_8_Index ? csrs_10_MAT : tlb_20_P0_MAT;
  wire [1:0] _GEN_1030 = 5'h15 == csrs_8_Index ? csrs_10_MAT : tlb_21_P0_MAT;
  wire [1:0] _GEN_1031 = 5'h16 == csrs_8_Index ? csrs_10_MAT : tlb_22_P0_MAT;
  wire [1:0] _GEN_1032 = 5'h17 == csrs_8_Index ? csrs_10_MAT : tlb_23_P0_MAT;
  wire [1:0] _GEN_1033 = 5'h18 == csrs_8_Index ? csrs_10_MAT : tlb_24_P0_MAT;
  wire [1:0] _GEN_1034 = 5'h19 == csrs_8_Index ? csrs_10_MAT : tlb_25_P0_MAT;
  wire [1:0] _GEN_1035 = 5'h1a == csrs_8_Index ? csrs_10_MAT : tlb_26_P0_MAT;
  wire [1:0] _GEN_1036 = 5'h1b == csrs_8_Index ? csrs_10_MAT : tlb_27_P0_MAT;
  wire [1:0] _GEN_1037 = 5'h1c == csrs_8_Index ? csrs_10_MAT : tlb_28_P0_MAT;
  wire [1:0] _GEN_1038 = 5'h1d == csrs_8_Index ? csrs_10_MAT : tlb_29_P0_MAT;
  wire [1:0] _GEN_1039 = 5'h1e == csrs_8_Index ? csrs_10_MAT : tlb_30_P0_MAT;
  wire [1:0] _GEN_1040 = 5'h1f == csrs_8_Index ? csrs_10_MAT : tlb_31_P0_MAT;
  wire  _GEN_1041 = 5'h0 == csrs_8_Index ? csrs_10_D : tlb_0_P0_D;
  wire  _GEN_1042 = 5'h1 == csrs_8_Index ? csrs_10_D : tlb_1_P0_D;
  wire  _GEN_1043 = 5'h2 == csrs_8_Index ? csrs_10_D : tlb_2_P0_D;
  wire  _GEN_1044 = 5'h3 == csrs_8_Index ? csrs_10_D : tlb_3_P0_D;
  wire  _GEN_1045 = 5'h4 == csrs_8_Index ? csrs_10_D : tlb_4_P0_D;
  wire  _GEN_1046 = 5'h5 == csrs_8_Index ? csrs_10_D : tlb_5_P0_D;
  wire  _GEN_1047 = 5'h6 == csrs_8_Index ? csrs_10_D : tlb_6_P0_D;
  wire  _GEN_1048 = 5'h7 == csrs_8_Index ? csrs_10_D : tlb_7_P0_D;
  wire  _GEN_1049 = 5'h8 == csrs_8_Index ? csrs_10_D : tlb_8_P0_D;
  wire  _GEN_1050 = 5'h9 == csrs_8_Index ? csrs_10_D : tlb_9_P0_D;
  wire  _GEN_1051 = 5'ha == csrs_8_Index ? csrs_10_D : tlb_10_P0_D;
  wire  _GEN_1052 = 5'hb == csrs_8_Index ? csrs_10_D : tlb_11_P0_D;
  wire  _GEN_1053 = 5'hc == csrs_8_Index ? csrs_10_D : tlb_12_P0_D;
  wire  _GEN_1054 = 5'hd == csrs_8_Index ? csrs_10_D : tlb_13_P0_D;
  wire  _GEN_1055 = 5'he == csrs_8_Index ? csrs_10_D : tlb_14_P0_D;
  wire  _GEN_1056 = 5'hf == csrs_8_Index ? csrs_10_D : tlb_15_P0_D;
  wire  _GEN_1057 = 5'h10 == csrs_8_Index ? csrs_10_D : tlb_16_P0_D;
  wire  _GEN_1058 = 5'h11 == csrs_8_Index ? csrs_10_D : tlb_17_P0_D;
  wire  _GEN_1059 = 5'h12 == csrs_8_Index ? csrs_10_D : tlb_18_P0_D;
  wire  _GEN_1060 = 5'h13 == csrs_8_Index ? csrs_10_D : tlb_19_P0_D;
  wire  _GEN_1061 = 5'h14 == csrs_8_Index ? csrs_10_D : tlb_20_P0_D;
  wire  _GEN_1062 = 5'h15 == csrs_8_Index ? csrs_10_D : tlb_21_P0_D;
  wire  _GEN_1063 = 5'h16 == csrs_8_Index ? csrs_10_D : tlb_22_P0_D;
  wire  _GEN_1064 = 5'h17 == csrs_8_Index ? csrs_10_D : tlb_23_P0_D;
  wire  _GEN_1065 = 5'h18 == csrs_8_Index ? csrs_10_D : tlb_24_P0_D;
  wire  _GEN_1066 = 5'h19 == csrs_8_Index ? csrs_10_D : tlb_25_P0_D;
  wire  _GEN_1067 = 5'h1a == csrs_8_Index ? csrs_10_D : tlb_26_P0_D;
  wire  _GEN_1068 = 5'h1b == csrs_8_Index ? csrs_10_D : tlb_27_P0_D;
  wire  _GEN_1069 = 5'h1c == csrs_8_Index ? csrs_10_D : tlb_28_P0_D;
  wire  _GEN_1070 = 5'h1d == csrs_8_Index ? csrs_10_D : tlb_29_P0_D;
  wire  _GEN_1071 = 5'h1e == csrs_8_Index ? csrs_10_D : tlb_30_P0_D;
  wire  _GEN_1072 = 5'h1f == csrs_8_Index ? csrs_10_D : tlb_31_P0_D;
  wire  _GEN_1073 = 5'h0 == csrs_8_Index ? csrs_10_V : tlb_0_P0_V;
  wire  _GEN_1074 = 5'h1 == csrs_8_Index ? csrs_10_V : tlb_1_P0_V;
  wire  _GEN_1075 = 5'h2 == csrs_8_Index ? csrs_10_V : tlb_2_P0_V;
  wire  _GEN_1076 = 5'h3 == csrs_8_Index ? csrs_10_V : tlb_3_P0_V;
  wire  _GEN_1077 = 5'h4 == csrs_8_Index ? csrs_10_V : tlb_4_P0_V;
  wire  _GEN_1078 = 5'h5 == csrs_8_Index ? csrs_10_V : tlb_5_P0_V;
  wire  _GEN_1079 = 5'h6 == csrs_8_Index ? csrs_10_V : tlb_6_P0_V;
  wire  _GEN_1080 = 5'h7 == csrs_8_Index ? csrs_10_V : tlb_7_P0_V;
  wire  _GEN_1081 = 5'h8 == csrs_8_Index ? csrs_10_V : tlb_8_P0_V;
  wire  _GEN_1082 = 5'h9 == csrs_8_Index ? csrs_10_V : tlb_9_P0_V;
  wire  _GEN_1083 = 5'ha == csrs_8_Index ? csrs_10_V : tlb_10_P0_V;
  wire  _GEN_1084 = 5'hb == csrs_8_Index ? csrs_10_V : tlb_11_P0_V;
  wire  _GEN_1085 = 5'hc == csrs_8_Index ? csrs_10_V : tlb_12_P0_V;
  wire  _GEN_1086 = 5'hd == csrs_8_Index ? csrs_10_V : tlb_13_P0_V;
  wire  _GEN_1087 = 5'he == csrs_8_Index ? csrs_10_V : tlb_14_P0_V;
  wire  _GEN_1088 = 5'hf == csrs_8_Index ? csrs_10_V : tlb_15_P0_V;
  wire  _GEN_1089 = 5'h10 == csrs_8_Index ? csrs_10_V : tlb_16_P0_V;
  wire  _GEN_1090 = 5'h11 == csrs_8_Index ? csrs_10_V : tlb_17_P0_V;
  wire  _GEN_1091 = 5'h12 == csrs_8_Index ? csrs_10_V : tlb_18_P0_V;
  wire  _GEN_1092 = 5'h13 == csrs_8_Index ? csrs_10_V : tlb_19_P0_V;
  wire  _GEN_1093 = 5'h14 == csrs_8_Index ? csrs_10_V : tlb_20_P0_V;
  wire  _GEN_1094 = 5'h15 == csrs_8_Index ? csrs_10_V : tlb_21_P0_V;
  wire  _GEN_1095 = 5'h16 == csrs_8_Index ? csrs_10_V : tlb_22_P0_V;
  wire  _GEN_1096 = 5'h17 == csrs_8_Index ? csrs_10_V : tlb_23_P0_V;
  wire  _GEN_1097 = 5'h18 == csrs_8_Index ? csrs_10_V : tlb_24_P0_V;
  wire  _GEN_1098 = 5'h19 == csrs_8_Index ? csrs_10_V : tlb_25_P0_V;
  wire  _GEN_1099 = 5'h1a == csrs_8_Index ? csrs_10_V : tlb_26_P0_V;
  wire  _GEN_1100 = 5'h1b == csrs_8_Index ? csrs_10_V : tlb_27_P0_V;
  wire  _GEN_1101 = 5'h1c == csrs_8_Index ? csrs_10_V : tlb_28_P0_V;
  wire  _GEN_1102 = 5'h1d == csrs_8_Index ? csrs_10_V : tlb_29_P0_V;
  wire  _GEN_1103 = 5'h1e == csrs_8_Index ? csrs_10_V : tlb_30_P0_V;
  wire  _GEN_1104 = 5'h1f == csrs_8_Index ? csrs_10_V : tlb_31_P0_V;
  wire [19:0] _GEN_1105 = 5'h0 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_0_P1_PPN;
  wire [19:0] _GEN_1106 = 5'h1 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_1_P1_PPN;
  wire [19:0] _GEN_1107 = 5'h2 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_2_P1_PPN;
  wire [19:0] _GEN_1108 = 5'h3 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_3_P1_PPN;
  wire [19:0] _GEN_1109 = 5'h4 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_4_P1_PPN;
  wire [19:0] _GEN_1110 = 5'h5 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_5_P1_PPN;
  wire [19:0] _GEN_1111 = 5'h6 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_6_P1_PPN;
  wire [19:0] _GEN_1112 = 5'h7 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_7_P1_PPN;
  wire [19:0] _GEN_1113 = 5'h8 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_8_P1_PPN;
  wire [19:0] _GEN_1114 = 5'h9 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_9_P1_PPN;
  wire [19:0] _GEN_1115 = 5'ha == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_10_P1_PPN;
  wire [19:0] _GEN_1116 = 5'hb == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_11_P1_PPN;
  wire [19:0] _GEN_1117 = 5'hc == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_12_P1_PPN;
  wire [19:0] _GEN_1118 = 5'hd == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_13_P1_PPN;
  wire [19:0] _GEN_1119 = 5'he == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_14_P1_PPN;
  wire [19:0] _GEN_1120 = 5'hf == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_15_P1_PPN;
  wire [19:0] _GEN_1121 = 5'h10 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_16_P1_PPN;
  wire [19:0] _GEN_1122 = 5'h11 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_17_P1_PPN;
  wire [19:0] _GEN_1123 = 5'h12 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_18_P1_PPN;
  wire [19:0] _GEN_1124 = 5'h13 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_19_P1_PPN;
  wire [19:0] _GEN_1125 = 5'h14 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_20_P1_PPN;
  wire [19:0] _GEN_1126 = 5'h15 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_21_P1_PPN;
  wire [19:0] _GEN_1127 = 5'h16 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_22_P1_PPN;
  wire [19:0] _GEN_1128 = 5'h17 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_23_P1_PPN;
  wire [19:0] _GEN_1129 = 5'h18 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_24_P1_PPN;
  wire [19:0] _GEN_1130 = 5'h19 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_25_P1_PPN;
  wire [19:0] _GEN_1131 = 5'h1a == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_26_P1_PPN;
  wire [19:0] _GEN_1132 = 5'h1b == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_27_P1_PPN;
  wire [19:0] _GEN_1133 = 5'h1c == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_28_P1_PPN;
  wire [19:0] _GEN_1134 = 5'h1d == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_29_P1_PPN;
  wire [19:0] _GEN_1135 = 5'h1e == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_30_P1_PPN;
  wire [19:0] _GEN_1136 = 5'h1f == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_31_P1_PPN;
  wire [1:0] _GEN_1137 = 5'h0 == csrs_8_Index ? csrs_11_PLV : tlb_0_P1_PLV;
  wire [1:0] _GEN_1138 = 5'h1 == csrs_8_Index ? csrs_11_PLV : tlb_1_P1_PLV;
  wire [1:0] _GEN_1139 = 5'h2 == csrs_8_Index ? csrs_11_PLV : tlb_2_P1_PLV;
  wire [1:0] _GEN_1140 = 5'h3 == csrs_8_Index ? csrs_11_PLV : tlb_3_P1_PLV;
  wire [1:0] _GEN_1141 = 5'h4 == csrs_8_Index ? csrs_11_PLV : tlb_4_P1_PLV;
  wire [1:0] _GEN_1142 = 5'h5 == csrs_8_Index ? csrs_11_PLV : tlb_5_P1_PLV;
  wire [1:0] _GEN_1143 = 5'h6 == csrs_8_Index ? csrs_11_PLV : tlb_6_P1_PLV;
  wire [1:0] _GEN_1144 = 5'h7 == csrs_8_Index ? csrs_11_PLV : tlb_7_P1_PLV;
  wire [1:0] _GEN_1145 = 5'h8 == csrs_8_Index ? csrs_11_PLV : tlb_8_P1_PLV;
  wire [1:0] _GEN_1146 = 5'h9 == csrs_8_Index ? csrs_11_PLV : tlb_9_P1_PLV;
  wire [1:0] _GEN_1147 = 5'ha == csrs_8_Index ? csrs_11_PLV : tlb_10_P1_PLV;
  wire [1:0] _GEN_1148 = 5'hb == csrs_8_Index ? csrs_11_PLV : tlb_11_P1_PLV;
  wire [1:0] _GEN_1149 = 5'hc == csrs_8_Index ? csrs_11_PLV : tlb_12_P1_PLV;
  wire [1:0] _GEN_1150 = 5'hd == csrs_8_Index ? csrs_11_PLV : tlb_13_P1_PLV;
  wire [1:0] _GEN_1151 = 5'he == csrs_8_Index ? csrs_11_PLV : tlb_14_P1_PLV;
  wire [1:0] _GEN_1152 = 5'hf == csrs_8_Index ? csrs_11_PLV : tlb_15_P1_PLV;
  wire [1:0] _GEN_1153 = 5'h10 == csrs_8_Index ? csrs_11_PLV : tlb_16_P1_PLV;
  wire [1:0] _GEN_1154 = 5'h11 == csrs_8_Index ? csrs_11_PLV : tlb_17_P1_PLV;
  wire [1:0] _GEN_1155 = 5'h12 == csrs_8_Index ? csrs_11_PLV : tlb_18_P1_PLV;
  wire [1:0] _GEN_1156 = 5'h13 == csrs_8_Index ? csrs_11_PLV : tlb_19_P1_PLV;
  wire [1:0] _GEN_1157 = 5'h14 == csrs_8_Index ? csrs_11_PLV : tlb_20_P1_PLV;
  wire [1:0] _GEN_1158 = 5'h15 == csrs_8_Index ? csrs_11_PLV : tlb_21_P1_PLV;
  wire [1:0] _GEN_1159 = 5'h16 == csrs_8_Index ? csrs_11_PLV : tlb_22_P1_PLV;
  wire [1:0] _GEN_1160 = 5'h17 == csrs_8_Index ? csrs_11_PLV : tlb_23_P1_PLV;
  wire [1:0] _GEN_1161 = 5'h18 == csrs_8_Index ? csrs_11_PLV : tlb_24_P1_PLV;
  wire [1:0] _GEN_1162 = 5'h19 == csrs_8_Index ? csrs_11_PLV : tlb_25_P1_PLV;
  wire [1:0] _GEN_1163 = 5'h1a == csrs_8_Index ? csrs_11_PLV : tlb_26_P1_PLV;
  wire [1:0] _GEN_1164 = 5'h1b == csrs_8_Index ? csrs_11_PLV : tlb_27_P1_PLV;
  wire [1:0] _GEN_1165 = 5'h1c == csrs_8_Index ? csrs_11_PLV : tlb_28_P1_PLV;
  wire [1:0] _GEN_1166 = 5'h1d == csrs_8_Index ? csrs_11_PLV : tlb_29_P1_PLV;
  wire [1:0] _GEN_1167 = 5'h1e == csrs_8_Index ? csrs_11_PLV : tlb_30_P1_PLV;
  wire [1:0] _GEN_1168 = 5'h1f == csrs_8_Index ? csrs_11_PLV : tlb_31_P1_PLV;
  wire [1:0] _GEN_1169 = 5'h0 == csrs_8_Index ? csrs_11_MAT : tlb_0_P1_MAT;
  wire [1:0] _GEN_1170 = 5'h1 == csrs_8_Index ? csrs_11_MAT : tlb_1_P1_MAT;
  wire [1:0] _GEN_1171 = 5'h2 == csrs_8_Index ? csrs_11_MAT : tlb_2_P1_MAT;
  wire [1:0] _GEN_1172 = 5'h3 == csrs_8_Index ? csrs_11_MAT : tlb_3_P1_MAT;
  wire [1:0] _GEN_1173 = 5'h4 == csrs_8_Index ? csrs_11_MAT : tlb_4_P1_MAT;
  wire [1:0] _GEN_1174 = 5'h5 == csrs_8_Index ? csrs_11_MAT : tlb_5_P1_MAT;
  wire [1:0] _GEN_1175 = 5'h6 == csrs_8_Index ? csrs_11_MAT : tlb_6_P1_MAT;
  wire [1:0] _GEN_1176 = 5'h7 == csrs_8_Index ? csrs_11_MAT : tlb_7_P1_MAT;
  wire [1:0] _GEN_1177 = 5'h8 == csrs_8_Index ? csrs_11_MAT : tlb_8_P1_MAT;
  wire [1:0] _GEN_1178 = 5'h9 == csrs_8_Index ? csrs_11_MAT : tlb_9_P1_MAT;
  wire [1:0] _GEN_1179 = 5'ha == csrs_8_Index ? csrs_11_MAT : tlb_10_P1_MAT;
  wire [1:0] _GEN_1180 = 5'hb == csrs_8_Index ? csrs_11_MAT : tlb_11_P1_MAT;
  wire [1:0] _GEN_1181 = 5'hc == csrs_8_Index ? csrs_11_MAT : tlb_12_P1_MAT;
  wire [1:0] _GEN_1182 = 5'hd == csrs_8_Index ? csrs_11_MAT : tlb_13_P1_MAT;
  wire [1:0] _GEN_1183 = 5'he == csrs_8_Index ? csrs_11_MAT : tlb_14_P1_MAT;
  wire [1:0] _GEN_1184 = 5'hf == csrs_8_Index ? csrs_11_MAT : tlb_15_P1_MAT;
  wire [1:0] _GEN_1185 = 5'h10 == csrs_8_Index ? csrs_11_MAT : tlb_16_P1_MAT;
  wire [1:0] _GEN_1186 = 5'h11 == csrs_8_Index ? csrs_11_MAT : tlb_17_P1_MAT;
  wire [1:0] _GEN_1187 = 5'h12 == csrs_8_Index ? csrs_11_MAT : tlb_18_P1_MAT;
  wire [1:0] _GEN_1188 = 5'h13 == csrs_8_Index ? csrs_11_MAT : tlb_19_P1_MAT;
  wire [1:0] _GEN_1189 = 5'h14 == csrs_8_Index ? csrs_11_MAT : tlb_20_P1_MAT;
  wire [1:0] _GEN_1190 = 5'h15 == csrs_8_Index ? csrs_11_MAT : tlb_21_P1_MAT;
  wire [1:0] _GEN_1191 = 5'h16 == csrs_8_Index ? csrs_11_MAT : tlb_22_P1_MAT;
  wire [1:0] _GEN_1192 = 5'h17 == csrs_8_Index ? csrs_11_MAT : tlb_23_P1_MAT;
  wire [1:0] _GEN_1193 = 5'h18 == csrs_8_Index ? csrs_11_MAT : tlb_24_P1_MAT;
  wire [1:0] _GEN_1194 = 5'h19 == csrs_8_Index ? csrs_11_MAT : tlb_25_P1_MAT;
  wire [1:0] _GEN_1195 = 5'h1a == csrs_8_Index ? csrs_11_MAT : tlb_26_P1_MAT;
  wire [1:0] _GEN_1196 = 5'h1b == csrs_8_Index ? csrs_11_MAT : tlb_27_P1_MAT;
  wire [1:0] _GEN_1197 = 5'h1c == csrs_8_Index ? csrs_11_MAT : tlb_28_P1_MAT;
  wire [1:0] _GEN_1198 = 5'h1d == csrs_8_Index ? csrs_11_MAT : tlb_29_P1_MAT;
  wire [1:0] _GEN_1199 = 5'h1e == csrs_8_Index ? csrs_11_MAT : tlb_30_P1_MAT;
  wire [1:0] _GEN_1200 = 5'h1f == csrs_8_Index ? csrs_11_MAT : tlb_31_P1_MAT;
  wire  _GEN_1201 = 5'h0 == csrs_8_Index ? csrs_11_D : tlb_0_P1_D;
  wire  _GEN_1202 = 5'h1 == csrs_8_Index ? csrs_11_D : tlb_1_P1_D;
  wire  _GEN_1203 = 5'h2 == csrs_8_Index ? csrs_11_D : tlb_2_P1_D;
  wire  _GEN_1204 = 5'h3 == csrs_8_Index ? csrs_11_D : tlb_3_P1_D;
  wire  _GEN_1205 = 5'h4 == csrs_8_Index ? csrs_11_D : tlb_4_P1_D;
  wire  _GEN_1206 = 5'h5 == csrs_8_Index ? csrs_11_D : tlb_5_P1_D;
  wire  _GEN_1207 = 5'h6 == csrs_8_Index ? csrs_11_D : tlb_6_P1_D;
  wire  _GEN_1208 = 5'h7 == csrs_8_Index ? csrs_11_D : tlb_7_P1_D;
  wire  _GEN_1209 = 5'h8 == csrs_8_Index ? csrs_11_D : tlb_8_P1_D;
  wire  _GEN_1210 = 5'h9 == csrs_8_Index ? csrs_11_D : tlb_9_P1_D;
  wire  _GEN_1211 = 5'ha == csrs_8_Index ? csrs_11_D : tlb_10_P1_D;
  wire  _GEN_1212 = 5'hb == csrs_8_Index ? csrs_11_D : tlb_11_P1_D;
  wire  _GEN_1213 = 5'hc == csrs_8_Index ? csrs_11_D : tlb_12_P1_D;
  wire  _GEN_1214 = 5'hd == csrs_8_Index ? csrs_11_D : tlb_13_P1_D;
  wire  _GEN_1215 = 5'he == csrs_8_Index ? csrs_11_D : tlb_14_P1_D;
  wire  _GEN_1216 = 5'hf == csrs_8_Index ? csrs_11_D : tlb_15_P1_D;
  wire  _GEN_1217 = 5'h10 == csrs_8_Index ? csrs_11_D : tlb_16_P1_D;
  wire  _GEN_1218 = 5'h11 == csrs_8_Index ? csrs_11_D : tlb_17_P1_D;
  wire  _GEN_1219 = 5'h12 == csrs_8_Index ? csrs_11_D : tlb_18_P1_D;
  wire  _GEN_1220 = 5'h13 == csrs_8_Index ? csrs_11_D : tlb_19_P1_D;
  wire  _GEN_1221 = 5'h14 == csrs_8_Index ? csrs_11_D : tlb_20_P1_D;
  wire  _GEN_1222 = 5'h15 == csrs_8_Index ? csrs_11_D : tlb_21_P1_D;
  wire  _GEN_1223 = 5'h16 == csrs_8_Index ? csrs_11_D : tlb_22_P1_D;
  wire  _GEN_1224 = 5'h17 == csrs_8_Index ? csrs_11_D : tlb_23_P1_D;
  wire  _GEN_1225 = 5'h18 == csrs_8_Index ? csrs_11_D : tlb_24_P1_D;
  wire  _GEN_1226 = 5'h19 == csrs_8_Index ? csrs_11_D : tlb_25_P1_D;
  wire  _GEN_1227 = 5'h1a == csrs_8_Index ? csrs_11_D : tlb_26_P1_D;
  wire  _GEN_1228 = 5'h1b == csrs_8_Index ? csrs_11_D : tlb_27_P1_D;
  wire  _GEN_1229 = 5'h1c == csrs_8_Index ? csrs_11_D : tlb_28_P1_D;
  wire  _GEN_1230 = 5'h1d == csrs_8_Index ? csrs_11_D : tlb_29_P1_D;
  wire  _GEN_1231 = 5'h1e == csrs_8_Index ? csrs_11_D : tlb_30_P1_D;
  wire  _GEN_1232 = 5'h1f == csrs_8_Index ? csrs_11_D : tlb_31_P1_D;
  wire  _GEN_1233 = 5'h0 == csrs_8_Index ? csrs_11_V : tlb_0_P1_V;
  wire  _GEN_1234 = 5'h1 == csrs_8_Index ? csrs_11_V : tlb_1_P1_V;
  wire  _GEN_1235 = 5'h2 == csrs_8_Index ? csrs_11_V : tlb_2_P1_V;
  wire  _GEN_1236 = 5'h3 == csrs_8_Index ? csrs_11_V : tlb_3_P1_V;
  wire  _GEN_1237 = 5'h4 == csrs_8_Index ? csrs_11_V : tlb_4_P1_V;
  wire  _GEN_1238 = 5'h5 == csrs_8_Index ? csrs_11_V : tlb_5_P1_V;
  wire  _GEN_1239 = 5'h6 == csrs_8_Index ? csrs_11_V : tlb_6_P1_V;
  wire  _GEN_1240 = 5'h7 == csrs_8_Index ? csrs_11_V : tlb_7_P1_V;
  wire  _GEN_1241 = 5'h8 == csrs_8_Index ? csrs_11_V : tlb_8_P1_V;
  wire  _GEN_1242 = 5'h9 == csrs_8_Index ? csrs_11_V : tlb_9_P1_V;
  wire  _GEN_1243 = 5'ha == csrs_8_Index ? csrs_11_V : tlb_10_P1_V;
  wire  _GEN_1244 = 5'hb == csrs_8_Index ? csrs_11_V : tlb_11_P1_V;
  wire  _GEN_1245 = 5'hc == csrs_8_Index ? csrs_11_V : tlb_12_P1_V;
  wire  _GEN_1246 = 5'hd == csrs_8_Index ? csrs_11_V : tlb_13_P1_V;
  wire  _GEN_1247 = 5'he == csrs_8_Index ? csrs_11_V : tlb_14_P1_V;
  wire  _GEN_1248 = 5'hf == csrs_8_Index ? csrs_11_V : tlb_15_P1_V;
  wire  _GEN_1249 = 5'h10 == csrs_8_Index ? csrs_11_V : tlb_16_P1_V;
  wire  _GEN_1250 = 5'h11 == csrs_8_Index ? csrs_11_V : tlb_17_P1_V;
  wire  _GEN_1251 = 5'h12 == csrs_8_Index ? csrs_11_V : tlb_18_P1_V;
  wire  _GEN_1252 = 5'h13 == csrs_8_Index ? csrs_11_V : tlb_19_P1_V;
  wire  _GEN_1253 = 5'h14 == csrs_8_Index ? csrs_11_V : tlb_20_P1_V;
  wire  _GEN_1254 = 5'h15 == csrs_8_Index ? csrs_11_V : tlb_21_P1_V;
  wire  _GEN_1255 = 5'h16 == csrs_8_Index ? csrs_11_V : tlb_22_P1_V;
  wire  _GEN_1256 = 5'h17 == csrs_8_Index ? csrs_11_V : tlb_23_P1_V;
  wire  _GEN_1257 = 5'h18 == csrs_8_Index ? csrs_11_V : tlb_24_P1_V;
  wire  _GEN_1258 = 5'h19 == csrs_8_Index ? csrs_11_V : tlb_25_P1_V;
  wire  _GEN_1259 = 5'h1a == csrs_8_Index ? csrs_11_V : tlb_26_P1_V;
  wire  _GEN_1260 = 5'h1b == csrs_8_Index ? csrs_11_V : tlb_27_P1_V;
  wire  _GEN_1261 = 5'h1c == csrs_8_Index ? csrs_11_V : tlb_28_P1_V;
  wire  _GEN_1262 = 5'h1d == csrs_8_Index ? csrs_11_V : tlb_29_P1_V;
  wire  _GEN_1263 = 5'h1e == csrs_8_Index ? csrs_11_V : tlb_30_P1_V;
  wire  _GEN_1264 = 5'h1f == csrs_8_Index ? csrs_11_V : tlb_31_P1_V;
  wire [18:0] _GEN_1265 = 5'h0 == timer[4:0] ? csrs_9_VPPN : tlb_0_VPPN;
  wire [18:0] _GEN_1266 = 5'h1 == timer[4:0] ? csrs_9_VPPN : tlb_1_VPPN;
  wire [18:0] _GEN_1267 = 5'h2 == timer[4:0] ? csrs_9_VPPN : tlb_2_VPPN;
  wire [18:0] _GEN_1268 = 5'h3 == timer[4:0] ? csrs_9_VPPN : tlb_3_VPPN;
  wire [18:0] _GEN_1269 = 5'h4 == timer[4:0] ? csrs_9_VPPN : tlb_4_VPPN;
  wire [18:0] _GEN_1270 = 5'h5 == timer[4:0] ? csrs_9_VPPN : tlb_5_VPPN;
  wire [18:0] _GEN_1271 = 5'h6 == timer[4:0] ? csrs_9_VPPN : tlb_6_VPPN;
  wire [18:0] _GEN_1272 = 5'h7 == timer[4:0] ? csrs_9_VPPN : tlb_7_VPPN;
  wire [18:0] _GEN_1273 = 5'h8 == timer[4:0] ? csrs_9_VPPN : tlb_8_VPPN;
  wire [18:0] _GEN_1274 = 5'h9 == timer[4:0] ? csrs_9_VPPN : tlb_9_VPPN;
  wire [18:0] _GEN_1275 = 5'ha == timer[4:0] ? csrs_9_VPPN : tlb_10_VPPN;
  wire [18:0] _GEN_1276 = 5'hb == timer[4:0] ? csrs_9_VPPN : tlb_11_VPPN;
  wire [18:0] _GEN_1277 = 5'hc == timer[4:0] ? csrs_9_VPPN : tlb_12_VPPN;
  wire [18:0] _GEN_1278 = 5'hd == timer[4:0] ? csrs_9_VPPN : tlb_13_VPPN;
  wire [18:0] _GEN_1279 = 5'he == timer[4:0] ? csrs_9_VPPN : tlb_14_VPPN;
  wire [18:0] _GEN_1280 = 5'hf == timer[4:0] ? csrs_9_VPPN : tlb_15_VPPN;
  wire [18:0] _GEN_1281 = 5'h10 == timer[4:0] ? csrs_9_VPPN : tlb_16_VPPN;
  wire [18:0] _GEN_1282 = 5'h11 == timer[4:0] ? csrs_9_VPPN : tlb_17_VPPN;
  wire [18:0] _GEN_1283 = 5'h12 == timer[4:0] ? csrs_9_VPPN : tlb_18_VPPN;
  wire [18:0] _GEN_1284 = 5'h13 == timer[4:0] ? csrs_9_VPPN : tlb_19_VPPN;
  wire [18:0] _GEN_1285 = 5'h14 == timer[4:0] ? csrs_9_VPPN : tlb_20_VPPN;
  wire [18:0] _GEN_1286 = 5'h15 == timer[4:0] ? csrs_9_VPPN : tlb_21_VPPN;
  wire [18:0] _GEN_1287 = 5'h16 == timer[4:0] ? csrs_9_VPPN : tlb_22_VPPN;
  wire [18:0] _GEN_1288 = 5'h17 == timer[4:0] ? csrs_9_VPPN : tlb_23_VPPN;
  wire [18:0] _GEN_1289 = 5'h18 == timer[4:0] ? csrs_9_VPPN : tlb_24_VPPN;
  wire [18:0] _GEN_1290 = 5'h19 == timer[4:0] ? csrs_9_VPPN : tlb_25_VPPN;
  wire [18:0] _GEN_1291 = 5'h1a == timer[4:0] ? csrs_9_VPPN : tlb_26_VPPN;
  wire [18:0] _GEN_1292 = 5'h1b == timer[4:0] ? csrs_9_VPPN : tlb_27_VPPN;
  wire [18:0] _GEN_1293 = 5'h1c == timer[4:0] ? csrs_9_VPPN : tlb_28_VPPN;
  wire [18:0] _GEN_1294 = 5'h1d == timer[4:0] ? csrs_9_VPPN : tlb_29_VPPN;
  wire [18:0] _GEN_1295 = 5'h1e == timer[4:0] ? csrs_9_VPPN : tlb_30_VPPN;
  wire [18:0] _GEN_1296 = 5'h1f == timer[4:0] ? csrs_9_VPPN : tlb_31_VPPN;
  wire [5:0] _GEN_1297 = 5'h0 == timer[4:0] ? csrs_8_PS : tlb_0_PS;
  wire [5:0] _GEN_1298 = 5'h1 == timer[4:0] ? csrs_8_PS : tlb_1_PS;
  wire [5:0] _GEN_1299 = 5'h2 == timer[4:0] ? csrs_8_PS : tlb_2_PS;
  wire [5:0] _GEN_1300 = 5'h3 == timer[4:0] ? csrs_8_PS : tlb_3_PS;
  wire [5:0] _GEN_1301 = 5'h4 == timer[4:0] ? csrs_8_PS : tlb_4_PS;
  wire [5:0] _GEN_1302 = 5'h5 == timer[4:0] ? csrs_8_PS : tlb_5_PS;
  wire [5:0] _GEN_1303 = 5'h6 == timer[4:0] ? csrs_8_PS : tlb_6_PS;
  wire [5:0] _GEN_1304 = 5'h7 == timer[4:0] ? csrs_8_PS : tlb_7_PS;
  wire [5:0] _GEN_1305 = 5'h8 == timer[4:0] ? csrs_8_PS : tlb_8_PS;
  wire [5:0] _GEN_1306 = 5'h9 == timer[4:0] ? csrs_8_PS : tlb_9_PS;
  wire [5:0] _GEN_1307 = 5'ha == timer[4:0] ? csrs_8_PS : tlb_10_PS;
  wire [5:0] _GEN_1308 = 5'hb == timer[4:0] ? csrs_8_PS : tlb_11_PS;
  wire [5:0] _GEN_1309 = 5'hc == timer[4:0] ? csrs_8_PS : tlb_12_PS;
  wire [5:0] _GEN_1310 = 5'hd == timer[4:0] ? csrs_8_PS : tlb_13_PS;
  wire [5:0] _GEN_1311 = 5'he == timer[4:0] ? csrs_8_PS : tlb_14_PS;
  wire [5:0] _GEN_1312 = 5'hf == timer[4:0] ? csrs_8_PS : tlb_15_PS;
  wire [5:0] _GEN_1313 = 5'h10 == timer[4:0] ? csrs_8_PS : tlb_16_PS;
  wire [5:0] _GEN_1314 = 5'h11 == timer[4:0] ? csrs_8_PS : tlb_17_PS;
  wire [5:0] _GEN_1315 = 5'h12 == timer[4:0] ? csrs_8_PS : tlb_18_PS;
  wire [5:0] _GEN_1316 = 5'h13 == timer[4:0] ? csrs_8_PS : tlb_19_PS;
  wire [5:0] _GEN_1317 = 5'h14 == timer[4:0] ? csrs_8_PS : tlb_20_PS;
  wire [5:0] _GEN_1318 = 5'h15 == timer[4:0] ? csrs_8_PS : tlb_21_PS;
  wire [5:0] _GEN_1319 = 5'h16 == timer[4:0] ? csrs_8_PS : tlb_22_PS;
  wire [5:0] _GEN_1320 = 5'h17 == timer[4:0] ? csrs_8_PS : tlb_23_PS;
  wire [5:0] _GEN_1321 = 5'h18 == timer[4:0] ? csrs_8_PS : tlb_24_PS;
  wire [5:0] _GEN_1322 = 5'h19 == timer[4:0] ? csrs_8_PS : tlb_25_PS;
  wire [5:0] _GEN_1323 = 5'h1a == timer[4:0] ? csrs_8_PS : tlb_26_PS;
  wire [5:0] _GEN_1324 = 5'h1b == timer[4:0] ? csrs_8_PS : tlb_27_PS;
  wire [5:0] _GEN_1325 = 5'h1c == timer[4:0] ? csrs_8_PS : tlb_28_PS;
  wire [5:0] _GEN_1326 = 5'h1d == timer[4:0] ? csrs_8_PS : tlb_29_PS;
  wire [5:0] _GEN_1327 = 5'h1e == timer[4:0] ? csrs_8_PS : tlb_30_PS;
  wire [5:0] _GEN_1328 = 5'h1f == timer[4:0] ? csrs_8_PS : tlb_31_PS;
  wire  _GEN_1329 = 5'h0 == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_0_G;
  wire  _GEN_1330 = 5'h1 == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_1_G;
  wire  _GEN_1331 = 5'h2 == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_2_G;
  wire  _GEN_1332 = 5'h3 == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_3_G;
  wire  _GEN_1333 = 5'h4 == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_4_G;
  wire  _GEN_1334 = 5'h5 == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_5_G;
  wire  _GEN_1335 = 5'h6 == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_6_G;
  wire  _GEN_1336 = 5'h7 == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_7_G;
  wire  _GEN_1337 = 5'h8 == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_8_G;
  wire  _GEN_1338 = 5'h9 == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_9_G;
  wire  _GEN_1339 = 5'ha == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_10_G;
  wire  _GEN_1340 = 5'hb == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_11_G;
  wire  _GEN_1341 = 5'hc == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_12_G;
  wire  _GEN_1342 = 5'hd == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_13_G;
  wire  _GEN_1343 = 5'he == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_14_G;
  wire  _GEN_1344 = 5'hf == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_15_G;
  wire  _GEN_1345 = 5'h10 == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_16_G;
  wire  _GEN_1346 = 5'h11 == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_17_G;
  wire  _GEN_1347 = 5'h12 == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_18_G;
  wire  _GEN_1348 = 5'h13 == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_19_G;
  wire  _GEN_1349 = 5'h14 == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_20_G;
  wire  _GEN_1350 = 5'h15 == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_21_G;
  wire  _GEN_1351 = 5'h16 == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_22_G;
  wire  _GEN_1352 = 5'h17 == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_23_G;
  wire  _GEN_1353 = 5'h18 == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_24_G;
  wire  _GEN_1354 = 5'h19 == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_25_G;
  wire  _GEN_1355 = 5'h1a == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_26_G;
  wire  _GEN_1356 = 5'h1b == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_27_G;
  wire  _GEN_1357 = 5'h1c == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_28_G;
  wire  _GEN_1358 = 5'h1d == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_29_G;
  wire  _GEN_1359 = 5'h1e == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_30_G;
  wire  _GEN_1360 = 5'h1f == timer[4:0] ? csrs_10_G & csrs_11_G : tlb_31_G;
  wire [9:0] _GEN_1361 = 5'h0 == timer[4:0] ? asid_ASID : tlb_0_ASID;
  wire [9:0] _GEN_1362 = 5'h1 == timer[4:0] ? asid_ASID : tlb_1_ASID;
  wire [9:0] _GEN_1363 = 5'h2 == timer[4:0] ? asid_ASID : tlb_2_ASID;
  wire [9:0] _GEN_1364 = 5'h3 == timer[4:0] ? asid_ASID : tlb_3_ASID;
  wire [9:0] _GEN_1365 = 5'h4 == timer[4:0] ? asid_ASID : tlb_4_ASID;
  wire [9:0] _GEN_1366 = 5'h5 == timer[4:0] ? asid_ASID : tlb_5_ASID;
  wire [9:0] _GEN_1367 = 5'h6 == timer[4:0] ? asid_ASID : tlb_6_ASID;
  wire [9:0] _GEN_1368 = 5'h7 == timer[4:0] ? asid_ASID : tlb_7_ASID;
  wire [9:0] _GEN_1369 = 5'h8 == timer[4:0] ? asid_ASID : tlb_8_ASID;
  wire [9:0] _GEN_1370 = 5'h9 == timer[4:0] ? asid_ASID : tlb_9_ASID;
  wire [9:0] _GEN_1371 = 5'ha == timer[4:0] ? asid_ASID : tlb_10_ASID;
  wire [9:0] _GEN_1372 = 5'hb == timer[4:0] ? asid_ASID : tlb_11_ASID;
  wire [9:0] _GEN_1373 = 5'hc == timer[4:0] ? asid_ASID : tlb_12_ASID;
  wire [9:0] _GEN_1374 = 5'hd == timer[4:0] ? asid_ASID : tlb_13_ASID;
  wire [9:0] _GEN_1375 = 5'he == timer[4:0] ? asid_ASID : tlb_14_ASID;
  wire [9:0] _GEN_1376 = 5'hf == timer[4:0] ? asid_ASID : tlb_15_ASID;
  wire [9:0] _GEN_1377 = 5'h10 == timer[4:0] ? asid_ASID : tlb_16_ASID;
  wire [9:0] _GEN_1378 = 5'h11 == timer[4:0] ? asid_ASID : tlb_17_ASID;
  wire [9:0] _GEN_1379 = 5'h12 == timer[4:0] ? asid_ASID : tlb_18_ASID;
  wire [9:0] _GEN_1380 = 5'h13 == timer[4:0] ? asid_ASID : tlb_19_ASID;
  wire [9:0] _GEN_1381 = 5'h14 == timer[4:0] ? asid_ASID : tlb_20_ASID;
  wire [9:0] _GEN_1382 = 5'h15 == timer[4:0] ? asid_ASID : tlb_21_ASID;
  wire [9:0] _GEN_1383 = 5'h16 == timer[4:0] ? asid_ASID : tlb_22_ASID;
  wire [9:0] _GEN_1384 = 5'h17 == timer[4:0] ? asid_ASID : tlb_23_ASID;
  wire [9:0] _GEN_1385 = 5'h18 == timer[4:0] ? asid_ASID : tlb_24_ASID;
  wire [9:0] _GEN_1386 = 5'h19 == timer[4:0] ? asid_ASID : tlb_25_ASID;
  wire [9:0] _GEN_1387 = 5'h1a == timer[4:0] ? asid_ASID : tlb_26_ASID;
  wire [9:0] _GEN_1388 = 5'h1b == timer[4:0] ? asid_ASID : tlb_27_ASID;
  wire [9:0] _GEN_1389 = 5'h1c == timer[4:0] ? asid_ASID : tlb_28_ASID;
  wire [9:0] _GEN_1390 = 5'h1d == timer[4:0] ? asid_ASID : tlb_29_ASID;
  wire [9:0] _GEN_1391 = 5'h1e == timer[4:0] ? asid_ASID : tlb_30_ASID;
  wire [9:0] _GEN_1392 = 5'h1f == timer[4:0] ? asid_ASID : tlb_31_ASID;
  wire  _GEN_1393 = 5'h0 == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_0_E;
  wire  _GEN_1394 = 5'h1 == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_1_E;
  wire  _GEN_1395 = 5'h2 == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_2_E;
  wire  _GEN_1396 = 5'h3 == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_3_E;
  wire  _GEN_1397 = 5'h4 == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_4_E;
  wire  _GEN_1398 = 5'h5 == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_5_E;
  wire  _GEN_1399 = 5'h6 == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_6_E;
  wire  _GEN_1400 = 5'h7 == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_7_E;
  wire  _GEN_1401 = 5'h8 == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_8_E;
  wire  _GEN_1402 = 5'h9 == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_9_E;
  wire  _GEN_1403 = 5'ha == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_10_E;
  wire  _GEN_1404 = 5'hb == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_11_E;
  wire  _GEN_1405 = 5'hc == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_12_E;
  wire  _GEN_1406 = 5'hd == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_13_E;
  wire  _GEN_1407 = 5'he == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_14_E;
  wire  _GEN_1408 = 5'hf == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_15_E;
  wire  _GEN_1409 = 5'h10 == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_16_E;
  wire  _GEN_1410 = 5'h11 == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_17_E;
  wire  _GEN_1411 = 5'h12 == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_18_E;
  wire  _GEN_1412 = 5'h13 == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_19_E;
  wire  _GEN_1413 = 5'h14 == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_20_E;
  wire  _GEN_1414 = 5'h15 == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_21_E;
  wire  _GEN_1415 = 5'h16 == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_22_E;
  wire  _GEN_1416 = 5'h17 == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_23_E;
  wire  _GEN_1417 = 5'h18 == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_24_E;
  wire  _GEN_1418 = 5'h19 == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_25_E;
  wire  _GEN_1419 = 5'h1a == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_26_E;
  wire  _GEN_1420 = 5'h1b == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_27_E;
  wire  _GEN_1421 = 5'h1c == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_28_E;
  wire  _GEN_1422 = 5'h1d == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_29_E;
  wire  _GEN_1423 = 5'h1e == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_30_E;
  wire  _GEN_1424 = 5'h1f == timer[4:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_31_E;
  wire [19:0] _GEN_1425 = 5'h0 == timer[4:0] ? csrs_10_PPN[19:0] : tlb_0_P0_PPN;
  wire [19:0] _GEN_1426 = 5'h1 == timer[4:0] ? csrs_10_PPN[19:0] : tlb_1_P0_PPN;
  wire [19:0] _GEN_1427 = 5'h2 == timer[4:0] ? csrs_10_PPN[19:0] : tlb_2_P0_PPN;
  wire [19:0] _GEN_1428 = 5'h3 == timer[4:0] ? csrs_10_PPN[19:0] : tlb_3_P0_PPN;
  wire [19:0] _GEN_1429 = 5'h4 == timer[4:0] ? csrs_10_PPN[19:0] : tlb_4_P0_PPN;
  wire [19:0] _GEN_1430 = 5'h5 == timer[4:0] ? csrs_10_PPN[19:0] : tlb_5_P0_PPN;
  wire [19:0] _GEN_1431 = 5'h6 == timer[4:0] ? csrs_10_PPN[19:0] : tlb_6_P0_PPN;
  wire [19:0] _GEN_1432 = 5'h7 == timer[4:0] ? csrs_10_PPN[19:0] : tlb_7_P0_PPN;
  wire [19:0] _GEN_1433 = 5'h8 == timer[4:0] ? csrs_10_PPN[19:0] : tlb_8_P0_PPN;
  wire [19:0] _GEN_1434 = 5'h9 == timer[4:0] ? csrs_10_PPN[19:0] : tlb_9_P0_PPN;
  wire [19:0] _GEN_1435 = 5'ha == timer[4:0] ? csrs_10_PPN[19:0] : tlb_10_P0_PPN;
  wire [19:0] _GEN_1436 = 5'hb == timer[4:0] ? csrs_10_PPN[19:0] : tlb_11_P0_PPN;
  wire [19:0] _GEN_1437 = 5'hc == timer[4:0] ? csrs_10_PPN[19:0] : tlb_12_P0_PPN;
  wire [19:0] _GEN_1438 = 5'hd == timer[4:0] ? csrs_10_PPN[19:0] : tlb_13_P0_PPN;
  wire [19:0] _GEN_1439 = 5'he == timer[4:0] ? csrs_10_PPN[19:0] : tlb_14_P0_PPN;
  wire [19:0] _GEN_1440 = 5'hf == timer[4:0] ? csrs_10_PPN[19:0] : tlb_15_P0_PPN;
  wire [19:0] _GEN_1441 = 5'h10 == timer[4:0] ? csrs_10_PPN[19:0] : tlb_16_P0_PPN;
  wire [19:0] _GEN_1442 = 5'h11 == timer[4:0] ? csrs_10_PPN[19:0] : tlb_17_P0_PPN;
  wire [19:0] _GEN_1443 = 5'h12 == timer[4:0] ? csrs_10_PPN[19:0] : tlb_18_P0_PPN;
  wire [19:0] _GEN_1444 = 5'h13 == timer[4:0] ? csrs_10_PPN[19:0] : tlb_19_P0_PPN;
  wire [19:0] _GEN_1445 = 5'h14 == timer[4:0] ? csrs_10_PPN[19:0] : tlb_20_P0_PPN;
  wire [19:0] _GEN_1446 = 5'h15 == timer[4:0] ? csrs_10_PPN[19:0] : tlb_21_P0_PPN;
  wire [19:0] _GEN_1447 = 5'h16 == timer[4:0] ? csrs_10_PPN[19:0] : tlb_22_P0_PPN;
  wire [19:0] _GEN_1448 = 5'h17 == timer[4:0] ? csrs_10_PPN[19:0] : tlb_23_P0_PPN;
  wire [19:0] _GEN_1449 = 5'h18 == timer[4:0] ? csrs_10_PPN[19:0] : tlb_24_P0_PPN;
  wire [19:0] _GEN_1450 = 5'h19 == timer[4:0] ? csrs_10_PPN[19:0] : tlb_25_P0_PPN;
  wire [19:0] _GEN_1451 = 5'h1a == timer[4:0] ? csrs_10_PPN[19:0] : tlb_26_P0_PPN;
  wire [19:0] _GEN_1452 = 5'h1b == timer[4:0] ? csrs_10_PPN[19:0] : tlb_27_P0_PPN;
  wire [19:0] _GEN_1453 = 5'h1c == timer[4:0] ? csrs_10_PPN[19:0] : tlb_28_P0_PPN;
  wire [19:0] _GEN_1454 = 5'h1d == timer[4:0] ? csrs_10_PPN[19:0] : tlb_29_P0_PPN;
  wire [19:0] _GEN_1455 = 5'h1e == timer[4:0] ? csrs_10_PPN[19:0] : tlb_30_P0_PPN;
  wire [19:0] _GEN_1456 = 5'h1f == timer[4:0] ? csrs_10_PPN[19:0] : tlb_31_P0_PPN;
  wire [1:0] _GEN_1457 = 5'h0 == timer[4:0] ? csrs_10_PLV : tlb_0_P0_PLV;
  wire [1:0] _GEN_1458 = 5'h1 == timer[4:0] ? csrs_10_PLV : tlb_1_P0_PLV;
  wire [1:0] _GEN_1459 = 5'h2 == timer[4:0] ? csrs_10_PLV : tlb_2_P0_PLV;
  wire [1:0] _GEN_1460 = 5'h3 == timer[4:0] ? csrs_10_PLV : tlb_3_P0_PLV;
  wire [1:0] _GEN_1461 = 5'h4 == timer[4:0] ? csrs_10_PLV : tlb_4_P0_PLV;
  wire [1:0] _GEN_1462 = 5'h5 == timer[4:0] ? csrs_10_PLV : tlb_5_P0_PLV;
  wire [1:0] _GEN_1463 = 5'h6 == timer[4:0] ? csrs_10_PLV : tlb_6_P0_PLV;
  wire [1:0] _GEN_1464 = 5'h7 == timer[4:0] ? csrs_10_PLV : tlb_7_P0_PLV;
  wire [1:0] _GEN_1465 = 5'h8 == timer[4:0] ? csrs_10_PLV : tlb_8_P0_PLV;
  wire [1:0] _GEN_1466 = 5'h9 == timer[4:0] ? csrs_10_PLV : tlb_9_P0_PLV;
  wire [1:0] _GEN_1467 = 5'ha == timer[4:0] ? csrs_10_PLV : tlb_10_P0_PLV;
  wire [1:0] _GEN_1468 = 5'hb == timer[4:0] ? csrs_10_PLV : tlb_11_P0_PLV;
  wire [1:0] _GEN_1469 = 5'hc == timer[4:0] ? csrs_10_PLV : tlb_12_P0_PLV;
  wire [1:0] _GEN_1470 = 5'hd == timer[4:0] ? csrs_10_PLV : tlb_13_P0_PLV;
  wire [1:0] _GEN_1471 = 5'he == timer[4:0] ? csrs_10_PLV : tlb_14_P0_PLV;
  wire [1:0] _GEN_1472 = 5'hf == timer[4:0] ? csrs_10_PLV : tlb_15_P0_PLV;
  wire [1:0] _GEN_1473 = 5'h10 == timer[4:0] ? csrs_10_PLV : tlb_16_P0_PLV;
  wire [1:0] _GEN_1474 = 5'h11 == timer[4:0] ? csrs_10_PLV : tlb_17_P0_PLV;
  wire [1:0] _GEN_1475 = 5'h12 == timer[4:0] ? csrs_10_PLV : tlb_18_P0_PLV;
  wire [1:0] _GEN_1476 = 5'h13 == timer[4:0] ? csrs_10_PLV : tlb_19_P0_PLV;
  wire [1:0] _GEN_1477 = 5'h14 == timer[4:0] ? csrs_10_PLV : tlb_20_P0_PLV;
  wire [1:0] _GEN_1478 = 5'h15 == timer[4:0] ? csrs_10_PLV : tlb_21_P0_PLV;
  wire [1:0] _GEN_1479 = 5'h16 == timer[4:0] ? csrs_10_PLV : tlb_22_P0_PLV;
  wire [1:0] _GEN_1480 = 5'h17 == timer[4:0] ? csrs_10_PLV : tlb_23_P0_PLV;
  wire [1:0] _GEN_1481 = 5'h18 == timer[4:0] ? csrs_10_PLV : tlb_24_P0_PLV;
  wire [1:0] _GEN_1482 = 5'h19 == timer[4:0] ? csrs_10_PLV : tlb_25_P0_PLV;
  wire [1:0] _GEN_1483 = 5'h1a == timer[4:0] ? csrs_10_PLV : tlb_26_P0_PLV;
  wire [1:0] _GEN_1484 = 5'h1b == timer[4:0] ? csrs_10_PLV : tlb_27_P0_PLV;
  wire [1:0] _GEN_1485 = 5'h1c == timer[4:0] ? csrs_10_PLV : tlb_28_P0_PLV;
  wire [1:0] _GEN_1486 = 5'h1d == timer[4:0] ? csrs_10_PLV : tlb_29_P0_PLV;
  wire [1:0] _GEN_1487 = 5'h1e == timer[4:0] ? csrs_10_PLV : tlb_30_P0_PLV;
  wire [1:0] _GEN_1488 = 5'h1f == timer[4:0] ? csrs_10_PLV : tlb_31_P0_PLV;
  wire [1:0] _GEN_1489 = 5'h0 == timer[4:0] ? csrs_10_MAT : tlb_0_P0_MAT;
  wire [1:0] _GEN_1490 = 5'h1 == timer[4:0] ? csrs_10_MAT : tlb_1_P0_MAT;
  wire [1:0] _GEN_1491 = 5'h2 == timer[4:0] ? csrs_10_MAT : tlb_2_P0_MAT;
  wire [1:0] _GEN_1492 = 5'h3 == timer[4:0] ? csrs_10_MAT : tlb_3_P0_MAT;
  wire [1:0] _GEN_1493 = 5'h4 == timer[4:0] ? csrs_10_MAT : tlb_4_P0_MAT;
  wire [1:0] _GEN_1494 = 5'h5 == timer[4:0] ? csrs_10_MAT : tlb_5_P0_MAT;
  wire [1:0] _GEN_1495 = 5'h6 == timer[4:0] ? csrs_10_MAT : tlb_6_P0_MAT;
  wire [1:0] _GEN_1496 = 5'h7 == timer[4:0] ? csrs_10_MAT : tlb_7_P0_MAT;
  wire [1:0] _GEN_1497 = 5'h8 == timer[4:0] ? csrs_10_MAT : tlb_8_P0_MAT;
  wire [1:0] _GEN_1498 = 5'h9 == timer[4:0] ? csrs_10_MAT : tlb_9_P0_MAT;
  wire [1:0] _GEN_1499 = 5'ha == timer[4:0] ? csrs_10_MAT : tlb_10_P0_MAT;
  wire [1:0] _GEN_1500 = 5'hb == timer[4:0] ? csrs_10_MAT : tlb_11_P0_MAT;
  wire [1:0] _GEN_1501 = 5'hc == timer[4:0] ? csrs_10_MAT : tlb_12_P0_MAT;
  wire [1:0] _GEN_1502 = 5'hd == timer[4:0] ? csrs_10_MAT : tlb_13_P0_MAT;
  wire [1:0] _GEN_1503 = 5'he == timer[4:0] ? csrs_10_MAT : tlb_14_P0_MAT;
  wire [1:0] _GEN_1504 = 5'hf == timer[4:0] ? csrs_10_MAT : tlb_15_P0_MAT;
  wire [1:0] _GEN_1505 = 5'h10 == timer[4:0] ? csrs_10_MAT : tlb_16_P0_MAT;
  wire [1:0] _GEN_1506 = 5'h11 == timer[4:0] ? csrs_10_MAT : tlb_17_P0_MAT;
  wire [1:0] _GEN_1507 = 5'h12 == timer[4:0] ? csrs_10_MAT : tlb_18_P0_MAT;
  wire [1:0] _GEN_1508 = 5'h13 == timer[4:0] ? csrs_10_MAT : tlb_19_P0_MAT;
  wire [1:0] _GEN_1509 = 5'h14 == timer[4:0] ? csrs_10_MAT : tlb_20_P0_MAT;
  wire [1:0] _GEN_1510 = 5'h15 == timer[4:0] ? csrs_10_MAT : tlb_21_P0_MAT;
  wire [1:0] _GEN_1511 = 5'h16 == timer[4:0] ? csrs_10_MAT : tlb_22_P0_MAT;
  wire [1:0] _GEN_1512 = 5'h17 == timer[4:0] ? csrs_10_MAT : tlb_23_P0_MAT;
  wire [1:0] _GEN_1513 = 5'h18 == timer[4:0] ? csrs_10_MAT : tlb_24_P0_MAT;
  wire [1:0] _GEN_1514 = 5'h19 == timer[4:0] ? csrs_10_MAT : tlb_25_P0_MAT;
  wire [1:0] _GEN_1515 = 5'h1a == timer[4:0] ? csrs_10_MAT : tlb_26_P0_MAT;
  wire [1:0] _GEN_1516 = 5'h1b == timer[4:0] ? csrs_10_MAT : tlb_27_P0_MAT;
  wire [1:0] _GEN_1517 = 5'h1c == timer[4:0] ? csrs_10_MAT : tlb_28_P0_MAT;
  wire [1:0] _GEN_1518 = 5'h1d == timer[4:0] ? csrs_10_MAT : tlb_29_P0_MAT;
  wire [1:0] _GEN_1519 = 5'h1e == timer[4:0] ? csrs_10_MAT : tlb_30_P0_MAT;
  wire [1:0] _GEN_1520 = 5'h1f == timer[4:0] ? csrs_10_MAT : tlb_31_P0_MAT;
  wire  _GEN_1521 = 5'h0 == timer[4:0] ? csrs_10_D : tlb_0_P0_D;
  wire  _GEN_1522 = 5'h1 == timer[4:0] ? csrs_10_D : tlb_1_P0_D;
  wire  _GEN_1523 = 5'h2 == timer[4:0] ? csrs_10_D : tlb_2_P0_D;
  wire  _GEN_1524 = 5'h3 == timer[4:0] ? csrs_10_D : tlb_3_P0_D;
  wire  _GEN_1525 = 5'h4 == timer[4:0] ? csrs_10_D : tlb_4_P0_D;
  wire  _GEN_1526 = 5'h5 == timer[4:0] ? csrs_10_D : tlb_5_P0_D;
  wire  _GEN_1527 = 5'h6 == timer[4:0] ? csrs_10_D : tlb_6_P0_D;
  wire  _GEN_1528 = 5'h7 == timer[4:0] ? csrs_10_D : tlb_7_P0_D;
  wire  _GEN_1529 = 5'h8 == timer[4:0] ? csrs_10_D : tlb_8_P0_D;
  wire  _GEN_1530 = 5'h9 == timer[4:0] ? csrs_10_D : tlb_9_P0_D;
  wire  _GEN_1531 = 5'ha == timer[4:0] ? csrs_10_D : tlb_10_P0_D;
  wire  _GEN_1532 = 5'hb == timer[4:0] ? csrs_10_D : tlb_11_P0_D;
  wire  _GEN_1533 = 5'hc == timer[4:0] ? csrs_10_D : tlb_12_P0_D;
  wire  _GEN_1534 = 5'hd == timer[4:0] ? csrs_10_D : tlb_13_P0_D;
  wire  _GEN_1535 = 5'he == timer[4:0] ? csrs_10_D : tlb_14_P0_D;
  wire  _GEN_1536 = 5'hf == timer[4:0] ? csrs_10_D : tlb_15_P0_D;
  wire  _GEN_1537 = 5'h10 == timer[4:0] ? csrs_10_D : tlb_16_P0_D;
  wire  _GEN_1538 = 5'h11 == timer[4:0] ? csrs_10_D : tlb_17_P0_D;
  wire  _GEN_1539 = 5'h12 == timer[4:0] ? csrs_10_D : tlb_18_P0_D;
  wire  _GEN_1540 = 5'h13 == timer[4:0] ? csrs_10_D : tlb_19_P0_D;
  wire  _GEN_1541 = 5'h14 == timer[4:0] ? csrs_10_D : tlb_20_P0_D;
  wire  _GEN_1542 = 5'h15 == timer[4:0] ? csrs_10_D : tlb_21_P0_D;
  wire  _GEN_1543 = 5'h16 == timer[4:0] ? csrs_10_D : tlb_22_P0_D;
  wire  _GEN_1544 = 5'h17 == timer[4:0] ? csrs_10_D : tlb_23_P0_D;
  wire  _GEN_1545 = 5'h18 == timer[4:0] ? csrs_10_D : tlb_24_P0_D;
  wire  _GEN_1546 = 5'h19 == timer[4:0] ? csrs_10_D : tlb_25_P0_D;
  wire  _GEN_1547 = 5'h1a == timer[4:0] ? csrs_10_D : tlb_26_P0_D;
  wire  _GEN_1548 = 5'h1b == timer[4:0] ? csrs_10_D : tlb_27_P0_D;
  wire  _GEN_1549 = 5'h1c == timer[4:0] ? csrs_10_D : tlb_28_P0_D;
  wire  _GEN_1550 = 5'h1d == timer[4:0] ? csrs_10_D : tlb_29_P0_D;
  wire  _GEN_1551 = 5'h1e == timer[4:0] ? csrs_10_D : tlb_30_P0_D;
  wire  _GEN_1552 = 5'h1f == timer[4:0] ? csrs_10_D : tlb_31_P0_D;
  wire  _GEN_1553 = 5'h0 == timer[4:0] ? csrs_10_V : tlb_0_P0_V;
  wire  _GEN_1554 = 5'h1 == timer[4:0] ? csrs_10_V : tlb_1_P0_V;
  wire  _GEN_1555 = 5'h2 == timer[4:0] ? csrs_10_V : tlb_2_P0_V;
  wire  _GEN_1556 = 5'h3 == timer[4:0] ? csrs_10_V : tlb_3_P0_V;
  wire  _GEN_1557 = 5'h4 == timer[4:0] ? csrs_10_V : tlb_4_P0_V;
  wire  _GEN_1558 = 5'h5 == timer[4:0] ? csrs_10_V : tlb_5_P0_V;
  wire  _GEN_1559 = 5'h6 == timer[4:0] ? csrs_10_V : tlb_6_P0_V;
  wire  _GEN_1560 = 5'h7 == timer[4:0] ? csrs_10_V : tlb_7_P0_V;
  wire  _GEN_1561 = 5'h8 == timer[4:0] ? csrs_10_V : tlb_8_P0_V;
  wire  _GEN_1562 = 5'h9 == timer[4:0] ? csrs_10_V : tlb_9_P0_V;
  wire  _GEN_1563 = 5'ha == timer[4:0] ? csrs_10_V : tlb_10_P0_V;
  wire  _GEN_1564 = 5'hb == timer[4:0] ? csrs_10_V : tlb_11_P0_V;
  wire  _GEN_1565 = 5'hc == timer[4:0] ? csrs_10_V : tlb_12_P0_V;
  wire  _GEN_1566 = 5'hd == timer[4:0] ? csrs_10_V : tlb_13_P0_V;
  wire  _GEN_1567 = 5'he == timer[4:0] ? csrs_10_V : tlb_14_P0_V;
  wire  _GEN_1568 = 5'hf == timer[4:0] ? csrs_10_V : tlb_15_P0_V;
  wire  _GEN_1569 = 5'h10 == timer[4:0] ? csrs_10_V : tlb_16_P0_V;
  wire  _GEN_1570 = 5'h11 == timer[4:0] ? csrs_10_V : tlb_17_P0_V;
  wire  _GEN_1571 = 5'h12 == timer[4:0] ? csrs_10_V : tlb_18_P0_V;
  wire  _GEN_1572 = 5'h13 == timer[4:0] ? csrs_10_V : tlb_19_P0_V;
  wire  _GEN_1573 = 5'h14 == timer[4:0] ? csrs_10_V : tlb_20_P0_V;
  wire  _GEN_1574 = 5'h15 == timer[4:0] ? csrs_10_V : tlb_21_P0_V;
  wire  _GEN_1575 = 5'h16 == timer[4:0] ? csrs_10_V : tlb_22_P0_V;
  wire  _GEN_1576 = 5'h17 == timer[4:0] ? csrs_10_V : tlb_23_P0_V;
  wire  _GEN_1577 = 5'h18 == timer[4:0] ? csrs_10_V : tlb_24_P0_V;
  wire  _GEN_1578 = 5'h19 == timer[4:0] ? csrs_10_V : tlb_25_P0_V;
  wire  _GEN_1579 = 5'h1a == timer[4:0] ? csrs_10_V : tlb_26_P0_V;
  wire  _GEN_1580 = 5'h1b == timer[4:0] ? csrs_10_V : tlb_27_P0_V;
  wire  _GEN_1581 = 5'h1c == timer[4:0] ? csrs_10_V : tlb_28_P0_V;
  wire  _GEN_1582 = 5'h1d == timer[4:0] ? csrs_10_V : tlb_29_P0_V;
  wire  _GEN_1583 = 5'h1e == timer[4:0] ? csrs_10_V : tlb_30_P0_V;
  wire  _GEN_1584 = 5'h1f == timer[4:0] ? csrs_10_V : tlb_31_P0_V;
  wire [19:0] _GEN_1585 = 5'h0 == timer[4:0] ? csrs_11_PPN[19:0] : tlb_0_P1_PPN;
  wire [19:0] _GEN_1586 = 5'h1 == timer[4:0] ? csrs_11_PPN[19:0] : tlb_1_P1_PPN;
  wire [19:0] _GEN_1587 = 5'h2 == timer[4:0] ? csrs_11_PPN[19:0] : tlb_2_P1_PPN;
  wire [19:0] _GEN_1588 = 5'h3 == timer[4:0] ? csrs_11_PPN[19:0] : tlb_3_P1_PPN;
  wire [19:0] _GEN_1589 = 5'h4 == timer[4:0] ? csrs_11_PPN[19:0] : tlb_4_P1_PPN;
  wire [19:0] _GEN_1590 = 5'h5 == timer[4:0] ? csrs_11_PPN[19:0] : tlb_5_P1_PPN;
  wire [19:0] _GEN_1591 = 5'h6 == timer[4:0] ? csrs_11_PPN[19:0] : tlb_6_P1_PPN;
  wire [19:0] _GEN_1592 = 5'h7 == timer[4:0] ? csrs_11_PPN[19:0] : tlb_7_P1_PPN;
  wire [19:0] _GEN_1593 = 5'h8 == timer[4:0] ? csrs_11_PPN[19:0] : tlb_8_P1_PPN;
  wire [19:0] _GEN_1594 = 5'h9 == timer[4:0] ? csrs_11_PPN[19:0] : tlb_9_P1_PPN;
  wire [19:0] _GEN_1595 = 5'ha == timer[4:0] ? csrs_11_PPN[19:0] : tlb_10_P1_PPN;
  wire [19:0] _GEN_1596 = 5'hb == timer[4:0] ? csrs_11_PPN[19:0] : tlb_11_P1_PPN;
  wire [19:0] _GEN_1597 = 5'hc == timer[4:0] ? csrs_11_PPN[19:0] : tlb_12_P1_PPN;
  wire [19:0] _GEN_1598 = 5'hd == timer[4:0] ? csrs_11_PPN[19:0] : tlb_13_P1_PPN;
  wire [19:0] _GEN_1599 = 5'he == timer[4:0] ? csrs_11_PPN[19:0] : tlb_14_P1_PPN;
  wire [19:0] _GEN_1600 = 5'hf == timer[4:0] ? csrs_11_PPN[19:0] : tlb_15_P1_PPN;
  wire [19:0] _GEN_1601 = 5'h10 == timer[4:0] ? csrs_11_PPN[19:0] : tlb_16_P1_PPN;
  wire [19:0] _GEN_1602 = 5'h11 == timer[4:0] ? csrs_11_PPN[19:0] : tlb_17_P1_PPN;
  wire [19:0] _GEN_1603 = 5'h12 == timer[4:0] ? csrs_11_PPN[19:0] : tlb_18_P1_PPN;
  wire [19:0] _GEN_1604 = 5'h13 == timer[4:0] ? csrs_11_PPN[19:0] : tlb_19_P1_PPN;
  wire [19:0] _GEN_1605 = 5'h14 == timer[4:0] ? csrs_11_PPN[19:0] : tlb_20_P1_PPN;
  wire [19:0] _GEN_1606 = 5'h15 == timer[4:0] ? csrs_11_PPN[19:0] : tlb_21_P1_PPN;
  wire [19:0] _GEN_1607 = 5'h16 == timer[4:0] ? csrs_11_PPN[19:0] : tlb_22_P1_PPN;
  wire [19:0] _GEN_1608 = 5'h17 == timer[4:0] ? csrs_11_PPN[19:0] : tlb_23_P1_PPN;
  wire [19:0] _GEN_1609 = 5'h18 == timer[4:0] ? csrs_11_PPN[19:0] : tlb_24_P1_PPN;
  wire [19:0] _GEN_1610 = 5'h19 == timer[4:0] ? csrs_11_PPN[19:0] : tlb_25_P1_PPN;
  wire [19:0] _GEN_1611 = 5'h1a == timer[4:0] ? csrs_11_PPN[19:0] : tlb_26_P1_PPN;
  wire [19:0] _GEN_1612 = 5'h1b == timer[4:0] ? csrs_11_PPN[19:0] : tlb_27_P1_PPN;
  wire [19:0] _GEN_1613 = 5'h1c == timer[4:0] ? csrs_11_PPN[19:0] : tlb_28_P1_PPN;
  wire [19:0] _GEN_1614 = 5'h1d == timer[4:0] ? csrs_11_PPN[19:0] : tlb_29_P1_PPN;
  wire [19:0] _GEN_1615 = 5'h1e == timer[4:0] ? csrs_11_PPN[19:0] : tlb_30_P1_PPN;
  wire [19:0] _GEN_1616 = 5'h1f == timer[4:0] ? csrs_11_PPN[19:0] : tlb_31_P1_PPN;
  wire [1:0] _GEN_1617 = 5'h0 == timer[4:0] ? csrs_11_PLV : tlb_0_P1_PLV;
  wire [1:0] _GEN_1618 = 5'h1 == timer[4:0] ? csrs_11_PLV : tlb_1_P1_PLV;
  wire [1:0] _GEN_1619 = 5'h2 == timer[4:0] ? csrs_11_PLV : tlb_2_P1_PLV;
  wire [1:0] _GEN_1620 = 5'h3 == timer[4:0] ? csrs_11_PLV : tlb_3_P1_PLV;
  wire [1:0] _GEN_1621 = 5'h4 == timer[4:0] ? csrs_11_PLV : tlb_4_P1_PLV;
  wire [1:0] _GEN_1622 = 5'h5 == timer[4:0] ? csrs_11_PLV : tlb_5_P1_PLV;
  wire [1:0] _GEN_1623 = 5'h6 == timer[4:0] ? csrs_11_PLV : tlb_6_P1_PLV;
  wire [1:0] _GEN_1624 = 5'h7 == timer[4:0] ? csrs_11_PLV : tlb_7_P1_PLV;
  wire [1:0] _GEN_1625 = 5'h8 == timer[4:0] ? csrs_11_PLV : tlb_8_P1_PLV;
  wire [1:0] _GEN_1626 = 5'h9 == timer[4:0] ? csrs_11_PLV : tlb_9_P1_PLV;
  wire [1:0] _GEN_1627 = 5'ha == timer[4:0] ? csrs_11_PLV : tlb_10_P1_PLV;
  wire [1:0] _GEN_1628 = 5'hb == timer[4:0] ? csrs_11_PLV : tlb_11_P1_PLV;
  wire [1:0] _GEN_1629 = 5'hc == timer[4:0] ? csrs_11_PLV : tlb_12_P1_PLV;
  wire [1:0] _GEN_1630 = 5'hd == timer[4:0] ? csrs_11_PLV : tlb_13_P1_PLV;
  wire [1:0] _GEN_1631 = 5'he == timer[4:0] ? csrs_11_PLV : tlb_14_P1_PLV;
  wire [1:0] _GEN_1632 = 5'hf == timer[4:0] ? csrs_11_PLV : tlb_15_P1_PLV;
  wire [1:0] _GEN_1633 = 5'h10 == timer[4:0] ? csrs_11_PLV : tlb_16_P1_PLV;
  wire [1:0] _GEN_1634 = 5'h11 == timer[4:0] ? csrs_11_PLV : tlb_17_P1_PLV;
  wire [1:0] _GEN_1635 = 5'h12 == timer[4:0] ? csrs_11_PLV : tlb_18_P1_PLV;
  wire [1:0] _GEN_1636 = 5'h13 == timer[4:0] ? csrs_11_PLV : tlb_19_P1_PLV;
  wire [1:0] _GEN_1637 = 5'h14 == timer[4:0] ? csrs_11_PLV : tlb_20_P1_PLV;
  wire [1:0] _GEN_1638 = 5'h15 == timer[4:0] ? csrs_11_PLV : tlb_21_P1_PLV;
  wire [1:0] _GEN_1639 = 5'h16 == timer[4:0] ? csrs_11_PLV : tlb_22_P1_PLV;
  wire [1:0] _GEN_1640 = 5'h17 == timer[4:0] ? csrs_11_PLV : tlb_23_P1_PLV;
  wire [1:0] _GEN_1641 = 5'h18 == timer[4:0] ? csrs_11_PLV : tlb_24_P1_PLV;
  wire [1:0] _GEN_1642 = 5'h19 == timer[4:0] ? csrs_11_PLV : tlb_25_P1_PLV;
  wire [1:0] _GEN_1643 = 5'h1a == timer[4:0] ? csrs_11_PLV : tlb_26_P1_PLV;
  wire [1:0] _GEN_1644 = 5'h1b == timer[4:0] ? csrs_11_PLV : tlb_27_P1_PLV;
  wire [1:0] _GEN_1645 = 5'h1c == timer[4:0] ? csrs_11_PLV : tlb_28_P1_PLV;
  wire [1:0] _GEN_1646 = 5'h1d == timer[4:0] ? csrs_11_PLV : tlb_29_P1_PLV;
  wire [1:0] _GEN_1647 = 5'h1e == timer[4:0] ? csrs_11_PLV : tlb_30_P1_PLV;
  wire [1:0] _GEN_1648 = 5'h1f == timer[4:0] ? csrs_11_PLV : tlb_31_P1_PLV;
  wire [1:0] _GEN_1649 = 5'h0 == timer[4:0] ? csrs_11_MAT : tlb_0_P1_MAT;
  wire [1:0] _GEN_1650 = 5'h1 == timer[4:0] ? csrs_11_MAT : tlb_1_P1_MAT;
  wire [1:0] _GEN_1651 = 5'h2 == timer[4:0] ? csrs_11_MAT : tlb_2_P1_MAT;
  wire [1:0] _GEN_1652 = 5'h3 == timer[4:0] ? csrs_11_MAT : tlb_3_P1_MAT;
  wire [1:0] _GEN_1653 = 5'h4 == timer[4:0] ? csrs_11_MAT : tlb_4_P1_MAT;
  wire [1:0] _GEN_1654 = 5'h5 == timer[4:0] ? csrs_11_MAT : tlb_5_P1_MAT;
  wire [1:0] _GEN_1655 = 5'h6 == timer[4:0] ? csrs_11_MAT : tlb_6_P1_MAT;
  wire [1:0] _GEN_1656 = 5'h7 == timer[4:0] ? csrs_11_MAT : tlb_7_P1_MAT;
  wire [1:0] _GEN_1657 = 5'h8 == timer[4:0] ? csrs_11_MAT : tlb_8_P1_MAT;
  wire [1:0] _GEN_1658 = 5'h9 == timer[4:0] ? csrs_11_MAT : tlb_9_P1_MAT;
  wire [1:0] _GEN_1659 = 5'ha == timer[4:0] ? csrs_11_MAT : tlb_10_P1_MAT;
  wire [1:0] _GEN_1660 = 5'hb == timer[4:0] ? csrs_11_MAT : tlb_11_P1_MAT;
  wire [1:0] _GEN_1661 = 5'hc == timer[4:0] ? csrs_11_MAT : tlb_12_P1_MAT;
  wire [1:0] _GEN_1662 = 5'hd == timer[4:0] ? csrs_11_MAT : tlb_13_P1_MAT;
  wire [1:0] _GEN_1663 = 5'he == timer[4:0] ? csrs_11_MAT : tlb_14_P1_MAT;
  wire [1:0] _GEN_1664 = 5'hf == timer[4:0] ? csrs_11_MAT : tlb_15_P1_MAT;
  wire [1:0] _GEN_1665 = 5'h10 == timer[4:0] ? csrs_11_MAT : tlb_16_P1_MAT;
  wire [1:0] _GEN_1666 = 5'h11 == timer[4:0] ? csrs_11_MAT : tlb_17_P1_MAT;
  wire [1:0] _GEN_1667 = 5'h12 == timer[4:0] ? csrs_11_MAT : tlb_18_P1_MAT;
  wire [1:0] _GEN_1668 = 5'h13 == timer[4:0] ? csrs_11_MAT : tlb_19_P1_MAT;
  wire [1:0] _GEN_1669 = 5'h14 == timer[4:0] ? csrs_11_MAT : tlb_20_P1_MAT;
  wire [1:0] _GEN_1670 = 5'h15 == timer[4:0] ? csrs_11_MAT : tlb_21_P1_MAT;
  wire [1:0] _GEN_1671 = 5'h16 == timer[4:0] ? csrs_11_MAT : tlb_22_P1_MAT;
  wire [1:0] _GEN_1672 = 5'h17 == timer[4:0] ? csrs_11_MAT : tlb_23_P1_MAT;
  wire [1:0] _GEN_1673 = 5'h18 == timer[4:0] ? csrs_11_MAT : tlb_24_P1_MAT;
  wire [1:0] _GEN_1674 = 5'h19 == timer[4:0] ? csrs_11_MAT : tlb_25_P1_MAT;
  wire [1:0] _GEN_1675 = 5'h1a == timer[4:0] ? csrs_11_MAT : tlb_26_P1_MAT;
  wire [1:0] _GEN_1676 = 5'h1b == timer[4:0] ? csrs_11_MAT : tlb_27_P1_MAT;
  wire [1:0] _GEN_1677 = 5'h1c == timer[4:0] ? csrs_11_MAT : tlb_28_P1_MAT;
  wire [1:0] _GEN_1678 = 5'h1d == timer[4:0] ? csrs_11_MAT : tlb_29_P1_MAT;
  wire [1:0] _GEN_1679 = 5'h1e == timer[4:0] ? csrs_11_MAT : tlb_30_P1_MAT;
  wire [1:0] _GEN_1680 = 5'h1f == timer[4:0] ? csrs_11_MAT : tlb_31_P1_MAT;
  wire  _GEN_1681 = 5'h0 == timer[4:0] ? csrs_11_D : tlb_0_P1_D;
  wire  _GEN_1682 = 5'h1 == timer[4:0] ? csrs_11_D : tlb_1_P1_D;
  wire  _GEN_1683 = 5'h2 == timer[4:0] ? csrs_11_D : tlb_2_P1_D;
  wire  _GEN_1684 = 5'h3 == timer[4:0] ? csrs_11_D : tlb_3_P1_D;
  wire  _GEN_1685 = 5'h4 == timer[4:0] ? csrs_11_D : tlb_4_P1_D;
  wire  _GEN_1686 = 5'h5 == timer[4:0] ? csrs_11_D : tlb_5_P1_D;
  wire  _GEN_1687 = 5'h6 == timer[4:0] ? csrs_11_D : tlb_6_P1_D;
  wire  _GEN_1688 = 5'h7 == timer[4:0] ? csrs_11_D : tlb_7_P1_D;
  wire  _GEN_1689 = 5'h8 == timer[4:0] ? csrs_11_D : tlb_8_P1_D;
  wire  _GEN_1690 = 5'h9 == timer[4:0] ? csrs_11_D : tlb_9_P1_D;
  wire  _GEN_1691 = 5'ha == timer[4:0] ? csrs_11_D : tlb_10_P1_D;
  wire  _GEN_1692 = 5'hb == timer[4:0] ? csrs_11_D : tlb_11_P1_D;
  wire  _GEN_1693 = 5'hc == timer[4:0] ? csrs_11_D : tlb_12_P1_D;
  wire  _GEN_1694 = 5'hd == timer[4:0] ? csrs_11_D : tlb_13_P1_D;
  wire  _GEN_1695 = 5'he == timer[4:0] ? csrs_11_D : tlb_14_P1_D;
  wire  _GEN_1696 = 5'hf == timer[4:0] ? csrs_11_D : tlb_15_P1_D;
  wire  _GEN_1697 = 5'h10 == timer[4:0] ? csrs_11_D : tlb_16_P1_D;
  wire  _GEN_1698 = 5'h11 == timer[4:0] ? csrs_11_D : tlb_17_P1_D;
  wire  _GEN_1699 = 5'h12 == timer[4:0] ? csrs_11_D : tlb_18_P1_D;
  wire  _GEN_1700 = 5'h13 == timer[4:0] ? csrs_11_D : tlb_19_P1_D;
  wire  _GEN_1701 = 5'h14 == timer[4:0] ? csrs_11_D : tlb_20_P1_D;
  wire  _GEN_1702 = 5'h15 == timer[4:0] ? csrs_11_D : tlb_21_P1_D;
  wire  _GEN_1703 = 5'h16 == timer[4:0] ? csrs_11_D : tlb_22_P1_D;
  wire  _GEN_1704 = 5'h17 == timer[4:0] ? csrs_11_D : tlb_23_P1_D;
  wire  _GEN_1705 = 5'h18 == timer[4:0] ? csrs_11_D : tlb_24_P1_D;
  wire  _GEN_1706 = 5'h19 == timer[4:0] ? csrs_11_D : tlb_25_P1_D;
  wire  _GEN_1707 = 5'h1a == timer[4:0] ? csrs_11_D : tlb_26_P1_D;
  wire  _GEN_1708 = 5'h1b == timer[4:0] ? csrs_11_D : tlb_27_P1_D;
  wire  _GEN_1709 = 5'h1c == timer[4:0] ? csrs_11_D : tlb_28_P1_D;
  wire  _GEN_1710 = 5'h1d == timer[4:0] ? csrs_11_D : tlb_29_P1_D;
  wire  _GEN_1711 = 5'h1e == timer[4:0] ? csrs_11_D : tlb_30_P1_D;
  wire  _GEN_1712 = 5'h1f == timer[4:0] ? csrs_11_D : tlb_31_P1_D;
  wire  _GEN_1713 = 5'h0 == timer[4:0] ? csrs_11_V : tlb_0_P1_V;
  wire  _GEN_1714 = 5'h1 == timer[4:0] ? csrs_11_V : tlb_1_P1_V;
  wire  _GEN_1715 = 5'h2 == timer[4:0] ? csrs_11_V : tlb_2_P1_V;
  wire  _GEN_1716 = 5'h3 == timer[4:0] ? csrs_11_V : tlb_3_P1_V;
  wire  _GEN_1717 = 5'h4 == timer[4:0] ? csrs_11_V : tlb_4_P1_V;
  wire  _GEN_1718 = 5'h5 == timer[4:0] ? csrs_11_V : tlb_5_P1_V;
  wire  _GEN_1719 = 5'h6 == timer[4:0] ? csrs_11_V : tlb_6_P1_V;
  wire  _GEN_1720 = 5'h7 == timer[4:0] ? csrs_11_V : tlb_7_P1_V;
  wire  _GEN_1721 = 5'h8 == timer[4:0] ? csrs_11_V : tlb_8_P1_V;
  wire  _GEN_1722 = 5'h9 == timer[4:0] ? csrs_11_V : tlb_9_P1_V;
  wire  _GEN_1723 = 5'ha == timer[4:0] ? csrs_11_V : tlb_10_P1_V;
  wire  _GEN_1724 = 5'hb == timer[4:0] ? csrs_11_V : tlb_11_P1_V;
  wire  _GEN_1725 = 5'hc == timer[4:0] ? csrs_11_V : tlb_12_P1_V;
  wire  _GEN_1726 = 5'hd == timer[4:0] ? csrs_11_V : tlb_13_P1_V;
  wire  _GEN_1727 = 5'he == timer[4:0] ? csrs_11_V : tlb_14_P1_V;
  wire  _GEN_1728 = 5'hf == timer[4:0] ? csrs_11_V : tlb_15_P1_V;
  wire  _GEN_1729 = 5'h10 == timer[4:0] ? csrs_11_V : tlb_16_P1_V;
  wire  _GEN_1730 = 5'h11 == timer[4:0] ? csrs_11_V : tlb_17_P1_V;
  wire  _GEN_1731 = 5'h12 == timer[4:0] ? csrs_11_V : tlb_18_P1_V;
  wire  _GEN_1732 = 5'h13 == timer[4:0] ? csrs_11_V : tlb_19_P1_V;
  wire  _GEN_1733 = 5'h14 == timer[4:0] ? csrs_11_V : tlb_20_P1_V;
  wire  _GEN_1734 = 5'h15 == timer[4:0] ? csrs_11_V : tlb_21_P1_V;
  wire  _GEN_1735 = 5'h16 == timer[4:0] ? csrs_11_V : tlb_22_P1_V;
  wire  _GEN_1736 = 5'h17 == timer[4:0] ? csrs_11_V : tlb_23_P1_V;
  wire  _GEN_1737 = 5'h18 == timer[4:0] ? csrs_11_V : tlb_24_P1_V;
  wire  _GEN_1738 = 5'h19 == timer[4:0] ? csrs_11_V : tlb_25_P1_V;
  wire  _GEN_1739 = 5'h1a == timer[4:0] ? csrs_11_V : tlb_26_P1_V;
  wire  _GEN_1740 = 5'h1b == timer[4:0] ? csrs_11_V : tlb_27_P1_V;
  wire  _GEN_1741 = 5'h1c == timer[4:0] ? csrs_11_V : tlb_28_P1_V;
  wire  _GEN_1742 = 5'h1d == timer[4:0] ? csrs_11_V : tlb_29_P1_V;
  wire  _GEN_1743 = 5'h1e == timer[4:0] ? csrs_11_V : tlb_30_P1_V;
  wire  _GEN_1744 = 5'h1f == timer[4:0] ? csrs_11_V : tlb_31_P1_V;
  wire  _tlb_0_E_T = ~tlb_0_G;
  wire  _tlb_0_E_T_2 = _tlb_0_E_T & asidMatch_0_1;
  wire  _tlb_0_E_T_5 = _tlb_0_E_T_2 & vaMatch_0_1;
  wire  _tlb_0_E_T_8 = (_tlb_0_E_T | asidMatch_0_1) & vaMatch_0_1;
  wire  _tlb_0_E_T_19 = inv_op_0 | inv_op_1 & tlb_0_G | inv_op_2 & _tlb_0_E_T | inv_op_3 & _tlb_0_E_T_2 | inv_op_4 &
    _tlb_0_E_T_5 | inv_op_5 & _tlb_0_E_T_8;
  wire  _tlb_1_E_T = ~tlb_1_G;
  wire  _tlb_1_E_T_2 = _tlb_1_E_T & asidMatch_1_1;
  wire  _tlb_1_E_T_5 = _tlb_1_E_T_2 & vaMatch_1_1;
  wire  _tlb_1_E_T_8 = (_tlb_1_E_T | asidMatch_1_1) & vaMatch_1_1;
  wire  _tlb_1_E_T_19 = inv_op_0 | inv_op_1 & tlb_1_G | inv_op_2 & _tlb_1_E_T | inv_op_3 & _tlb_1_E_T_2 | inv_op_4 &
    _tlb_1_E_T_5 | inv_op_5 & _tlb_1_E_T_8;
  wire  _tlb_2_E_T = ~tlb_2_G;
  wire  _tlb_2_E_T_2 = _tlb_2_E_T & asidMatch_2_1;
  wire  _tlb_2_E_T_5 = _tlb_2_E_T_2 & vaMatch_2_1;
  wire  _tlb_2_E_T_8 = (_tlb_2_E_T | asidMatch_2_1) & vaMatch_2_1;
  wire  _tlb_2_E_T_19 = inv_op_0 | inv_op_1 & tlb_2_G | inv_op_2 & _tlb_2_E_T | inv_op_3 & _tlb_2_E_T_2 | inv_op_4 &
    _tlb_2_E_T_5 | inv_op_5 & _tlb_2_E_T_8;
  wire  _tlb_3_E_T = ~tlb_3_G;
  wire  _tlb_3_E_T_2 = _tlb_3_E_T & asidMatch_3_1;
  wire  _tlb_3_E_T_5 = _tlb_3_E_T_2 & vaMatch_3_1;
  wire  _tlb_3_E_T_8 = (_tlb_3_E_T | asidMatch_3_1) & vaMatch_3_1;
  wire  _tlb_3_E_T_19 = inv_op_0 | inv_op_1 & tlb_3_G | inv_op_2 & _tlb_3_E_T | inv_op_3 & _tlb_3_E_T_2 | inv_op_4 &
    _tlb_3_E_T_5 | inv_op_5 & _tlb_3_E_T_8;
  wire  _tlb_4_E_T = ~tlb_4_G;
  wire  _tlb_4_E_T_2 = _tlb_4_E_T & asidMatch_4_1;
  wire  _tlb_4_E_T_5 = _tlb_4_E_T_2 & vaMatch_4_1;
  wire  _tlb_4_E_T_8 = (_tlb_4_E_T | asidMatch_4_1) & vaMatch_4_1;
  wire  _tlb_4_E_T_19 = inv_op_0 | inv_op_1 & tlb_4_G | inv_op_2 & _tlb_4_E_T | inv_op_3 & _tlb_4_E_T_2 | inv_op_4 &
    _tlb_4_E_T_5 | inv_op_5 & _tlb_4_E_T_8;
  wire  _tlb_5_E_T = ~tlb_5_G;
  wire  _tlb_5_E_T_2 = _tlb_5_E_T & asidMatch_5_1;
  wire  _tlb_5_E_T_5 = _tlb_5_E_T_2 & vaMatch_5_1;
  wire  _tlb_5_E_T_8 = (_tlb_5_E_T | asidMatch_5_1) & vaMatch_5_1;
  wire  _tlb_5_E_T_19 = inv_op_0 | inv_op_1 & tlb_5_G | inv_op_2 & _tlb_5_E_T | inv_op_3 & _tlb_5_E_T_2 | inv_op_4 &
    _tlb_5_E_T_5 | inv_op_5 & _tlb_5_E_T_8;
  wire  _tlb_6_E_T = ~tlb_6_G;
  wire  _tlb_6_E_T_2 = _tlb_6_E_T & asidMatch_6_1;
  wire  _tlb_6_E_T_5 = _tlb_6_E_T_2 & vaMatch_6_1;
  wire  _tlb_6_E_T_8 = (_tlb_6_E_T | asidMatch_6_1) & vaMatch_6_1;
  wire  _tlb_6_E_T_19 = inv_op_0 | inv_op_1 & tlb_6_G | inv_op_2 & _tlb_6_E_T | inv_op_3 & _tlb_6_E_T_2 | inv_op_4 &
    _tlb_6_E_T_5 | inv_op_5 & _tlb_6_E_T_8;
  wire  _tlb_7_E_T = ~tlb_7_G;
  wire  _tlb_7_E_T_2 = _tlb_7_E_T & asidMatch_7_1;
  wire  _tlb_7_E_T_5 = _tlb_7_E_T_2 & vaMatch_7_1;
  wire  _tlb_7_E_T_8 = (_tlb_7_E_T | asidMatch_7_1) & vaMatch_7_1;
  wire  _tlb_7_E_T_19 = inv_op_0 | inv_op_1 & tlb_7_G | inv_op_2 & _tlb_7_E_T | inv_op_3 & _tlb_7_E_T_2 | inv_op_4 &
    _tlb_7_E_T_5 | inv_op_5 & _tlb_7_E_T_8;
  wire  _tlb_8_E_T = ~tlb_8_G;
  wire  _tlb_8_E_T_2 = _tlb_8_E_T & asidMatch_8_1;
  wire  _tlb_8_E_T_5 = _tlb_8_E_T_2 & vaMatch_8_1;
  wire  _tlb_8_E_T_8 = (_tlb_8_E_T | asidMatch_8_1) & vaMatch_8_1;
  wire  _tlb_8_E_T_19 = inv_op_0 | inv_op_1 & tlb_8_G | inv_op_2 & _tlb_8_E_T | inv_op_3 & _tlb_8_E_T_2 | inv_op_4 &
    _tlb_8_E_T_5 | inv_op_5 & _tlb_8_E_T_8;
  wire  _tlb_9_E_T = ~tlb_9_G;
  wire  _tlb_9_E_T_2 = _tlb_9_E_T & asidMatch_9_1;
  wire  _tlb_9_E_T_5 = _tlb_9_E_T_2 & vaMatch_9_1;
  wire  _tlb_9_E_T_8 = (_tlb_9_E_T | asidMatch_9_1) & vaMatch_9_1;
  wire  _tlb_9_E_T_19 = inv_op_0 | inv_op_1 & tlb_9_G | inv_op_2 & _tlb_9_E_T | inv_op_3 & _tlb_9_E_T_2 | inv_op_4 &
    _tlb_9_E_T_5 | inv_op_5 & _tlb_9_E_T_8;
  wire  _tlb_10_E_T = ~tlb_10_G;
  wire  _tlb_10_E_T_2 = _tlb_10_E_T & asidMatch_10_1;
  wire  _tlb_10_E_T_5 = _tlb_10_E_T_2 & vaMatch_10_1;
  wire  _tlb_10_E_T_8 = (_tlb_10_E_T | asidMatch_10_1) & vaMatch_10_1;
  wire  _tlb_10_E_T_19 = inv_op_0 | inv_op_1 & tlb_10_G | inv_op_2 & _tlb_10_E_T | inv_op_3 & _tlb_10_E_T_2 | inv_op_4
     & _tlb_10_E_T_5 | inv_op_5 & _tlb_10_E_T_8;
  wire  _tlb_11_E_T = ~tlb_11_G;
  wire  _tlb_11_E_T_2 = _tlb_11_E_T & asidMatch_11_1;
  wire  _tlb_11_E_T_5 = _tlb_11_E_T_2 & vaMatch_11_1;
  wire  _tlb_11_E_T_8 = (_tlb_11_E_T | asidMatch_11_1) & vaMatch_11_1;
  wire  _tlb_11_E_T_19 = inv_op_0 | inv_op_1 & tlb_11_G | inv_op_2 & _tlb_11_E_T | inv_op_3 & _tlb_11_E_T_2 | inv_op_4
     & _tlb_11_E_T_5 | inv_op_5 & _tlb_11_E_T_8;
  wire  _tlb_12_E_T = ~tlb_12_G;
  wire  _tlb_12_E_T_2 = _tlb_12_E_T & asidMatch_12_1;
  wire  _tlb_12_E_T_5 = _tlb_12_E_T_2 & vaMatch_12_1;
  wire  _tlb_12_E_T_8 = (_tlb_12_E_T | asidMatch_12_1) & vaMatch_12_1;
  wire  _tlb_12_E_T_19 = inv_op_0 | inv_op_1 & tlb_12_G | inv_op_2 & _tlb_12_E_T | inv_op_3 & _tlb_12_E_T_2 | inv_op_4
     & _tlb_12_E_T_5 | inv_op_5 & _tlb_12_E_T_8;
  wire  _tlb_13_E_T = ~tlb_13_G;
  wire  _tlb_13_E_T_2 = _tlb_13_E_T & asidMatch_13_1;
  wire  _tlb_13_E_T_5 = _tlb_13_E_T_2 & vaMatch_13_1;
  wire  _tlb_13_E_T_8 = (_tlb_13_E_T | asidMatch_13_1) & vaMatch_13_1;
  wire  _tlb_13_E_T_19 = inv_op_0 | inv_op_1 & tlb_13_G | inv_op_2 & _tlb_13_E_T | inv_op_3 & _tlb_13_E_T_2 | inv_op_4
     & _tlb_13_E_T_5 | inv_op_5 & _tlb_13_E_T_8;
  wire  _tlb_14_E_T = ~tlb_14_G;
  wire  _tlb_14_E_T_2 = _tlb_14_E_T & asidMatch_14_1;
  wire  _tlb_14_E_T_5 = _tlb_14_E_T_2 & vaMatch_14_1;
  wire  _tlb_14_E_T_8 = (_tlb_14_E_T | asidMatch_14_1) & vaMatch_14_1;
  wire  _tlb_14_E_T_19 = inv_op_0 | inv_op_1 & tlb_14_G | inv_op_2 & _tlb_14_E_T | inv_op_3 & _tlb_14_E_T_2 | inv_op_4
     & _tlb_14_E_T_5 | inv_op_5 & _tlb_14_E_T_8;
  wire  _tlb_15_E_T = ~tlb_15_G;
  wire  _tlb_15_E_T_2 = _tlb_15_E_T & asidMatch_15_1;
  wire  _tlb_15_E_T_5 = _tlb_15_E_T_2 & vaMatch_15_1;
  wire  _tlb_15_E_T_8 = (_tlb_15_E_T | asidMatch_15_1) & vaMatch_15_1;
  wire  _tlb_15_E_T_19 = inv_op_0 | inv_op_1 & tlb_15_G | inv_op_2 & _tlb_15_E_T | inv_op_3 & _tlb_15_E_T_2 | inv_op_4
     & _tlb_15_E_T_5 | inv_op_5 & _tlb_15_E_T_8;
  wire  _tlb_16_E_T = ~tlb_16_G;
  wire  _tlb_16_E_T_2 = _tlb_16_E_T & asidMatch_16_1;
  wire  _tlb_16_E_T_5 = _tlb_16_E_T_2 & vaMatch_16_1;
  wire  _tlb_16_E_T_8 = (_tlb_16_E_T | asidMatch_16_1) & vaMatch_16_1;
  wire  _tlb_16_E_T_19 = inv_op_0 | inv_op_1 & tlb_16_G | inv_op_2 & _tlb_16_E_T | inv_op_3 & _tlb_16_E_T_2 | inv_op_4
     & _tlb_16_E_T_5 | inv_op_5 & _tlb_16_E_T_8;
  wire  _tlb_17_E_T = ~tlb_17_G;
  wire  _tlb_17_E_T_2 = _tlb_17_E_T & asidMatch_17_1;
  wire  _tlb_17_E_T_5 = _tlb_17_E_T_2 & vaMatch_17_1;
  wire  _tlb_17_E_T_8 = (_tlb_17_E_T | asidMatch_17_1) & vaMatch_17_1;
  wire  _tlb_17_E_T_19 = inv_op_0 | inv_op_1 & tlb_17_G | inv_op_2 & _tlb_17_E_T | inv_op_3 & _tlb_17_E_T_2 | inv_op_4
     & _tlb_17_E_T_5 | inv_op_5 & _tlb_17_E_T_8;
  wire  _tlb_18_E_T = ~tlb_18_G;
  wire  _tlb_18_E_T_2 = _tlb_18_E_T & asidMatch_18_1;
  wire  _tlb_18_E_T_5 = _tlb_18_E_T_2 & vaMatch_18_1;
  wire  _tlb_18_E_T_8 = (_tlb_18_E_T | asidMatch_18_1) & vaMatch_18_1;
  wire  _tlb_18_E_T_19 = inv_op_0 | inv_op_1 & tlb_18_G | inv_op_2 & _tlb_18_E_T | inv_op_3 & _tlb_18_E_T_2 | inv_op_4
     & _tlb_18_E_T_5 | inv_op_5 & _tlb_18_E_T_8;
  wire  _tlb_19_E_T = ~tlb_19_G;
  wire  _tlb_19_E_T_2 = _tlb_19_E_T & asidMatch_19_1;
  wire  _tlb_19_E_T_5 = _tlb_19_E_T_2 & vaMatch_19_1;
  wire  _tlb_19_E_T_8 = (_tlb_19_E_T | asidMatch_19_1) & vaMatch_19_1;
  wire  _tlb_19_E_T_19 = inv_op_0 | inv_op_1 & tlb_19_G | inv_op_2 & _tlb_19_E_T | inv_op_3 & _tlb_19_E_T_2 | inv_op_4
     & _tlb_19_E_T_5 | inv_op_5 & _tlb_19_E_T_8;
  wire  _tlb_20_E_T = ~tlb_20_G;
  wire  _tlb_20_E_T_2 = _tlb_20_E_T & asidMatch_20_1;
  wire  _tlb_20_E_T_5 = _tlb_20_E_T_2 & vaMatch_20_1;
  wire  _tlb_20_E_T_8 = (_tlb_20_E_T | asidMatch_20_1) & vaMatch_20_1;
  wire  _tlb_20_E_T_19 = inv_op_0 | inv_op_1 & tlb_20_G | inv_op_2 & _tlb_20_E_T | inv_op_3 & _tlb_20_E_T_2 | inv_op_4
     & _tlb_20_E_T_5 | inv_op_5 & _tlb_20_E_T_8;
  wire  _tlb_21_E_T = ~tlb_21_G;
  wire  _tlb_21_E_T_2 = _tlb_21_E_T & asidMatch_21_1;
  wire  _tlb_21_E_T_5 = _tlb_21_E_T_2 & vaMatch_21_1;
  wire  _tlb_21_E_T_8 = (_tlb_21_E_T | asidMatch_21_1) & vaMatch_21_1;
  wire  _tlb_21_E_T_19 = inv_op_0 | inv_op_1 & tlb_21_G | inv_op_2 & _tlb_21_E_T | inv_op_3 & _tlb_21_E_T_2 | inv_op_4
     & _tlb_21_E_T_5 | inv_op_5 & _tlb_21_E_T_8;
  wire  _tlb_22_E_T = ~tlb_22_G;
  wire  _tlb_22_E_T_2 = _tlb_22_E_T & asidMatch_22_1;
  wire  _tlb_22_E_T_5 = _tlb_22_E_T_2 & vaMatch_22_1;
  wire  _tlb_22_E_T_8 = (_tlb_22_E_T | asidMatch_22_1) & vaMatch_22_1;
  wire  _tlb_22_E_T_19 = inv_op_0 | inv_op_1 & tlb_22_G | inv_op_2 & _tlb_22_E_T | inv_op_3 & _tlb_22_E_T_2 | inv_op_4
     & _tlb_22_E_T_5 | inv_op_5 & _tlb_22_E_T_8;
  wire  _tlb_23_E_T = ~tlb_23_G;
  wire  _tlb_23_E_T_2 = _tlb_23_E_T & asidMatch_23_1;
  wire  _tlb_23_E_T_5 = _tlb_23_E_T_2 & vaMatch_23_1;
  wire  _tlb_23_E_T_8 = (_tlb_23_E_T | asidMatch_23_1) & vaMatch_23_1;
  wire  _tlb_23_E_T_19 = inv_op_0 | inv_op_1 & tlb_23_G | inv_op_2 & _tlb_23_E_T | inv_op_3 & _tlb_23_E_T_2 | inv_op_4
     & _tlb_23_E_T_5 | inv_op_5 & _tlb_23_E_T_8;
  wire  _tlb_24_E_T = ~tlb_24_G;
  wire  _tlb_24_E_T_2 = _tlb_24_E_T & asidMatch_24_1;
  wire  _tlb_24_E_T_5 = _tlb_24_E_T_2 & vaMatch_24_1;
  wire  _tlb_24_E_T_8 = (_tlb_24_E_T | asidMatch_24_1) & vaMatch_24_1;
  wire  _tlb_24_E_T_19 = inv_op_0 | inv_op_1 & tlb_24_G | inv_op_2 & _tlb_24_E_T | inv_op_3 & _tlb_24_E_T_2 | inv_op_4
     & _tlb_24_E_T_5 | inv_op_5 & _tlb_24_E_T_8;
  wire  _tlb_25_E_T = ~tlb_25_G;
  wire  _tlb_25_E_T_2 = _tlb_25_E_T & asidMatch_25_1;
  wire  _tlb_25_E_T_5 = _tlb_25_E_T_2 & vaMatch_25_1;
  wire  _tlb_25_E_T_8 = (_tlb_25_E_T | asidMatch_25_1) & vaMatch_25_1;
  wire  _tlb_25_E_T_19 = inv_op_0 | inv_op_1 & tlb_25_G | inv_op_2 & _tlb_25_E_T | inv_op_3 & _tlb_25_E_T_2 | inv_op_4
     & _tlb_25_E_T_5 | inv_op_5 & _tlb_25_E_T_8;
  wire  _tlb_26_E_T = ~tlb_26_G;
  wire  _tlb_26_E_T_2 = _tlb_26_E_T & asidMatch_26_1;
  wire  _tlb_26_E_T_5 = _tlb_26_E_T_2 & vaMatch_26_1;
  wire  _tlb_26_E_T_8 = (_tlb_26_E_T | asidMatch_26_1) & vaMatch_26_1;
  wire  _tlb_26_E_T_19 = inv_op_0 | inv_op_1 & tlb_26_G | inv_op_2 & _tlb_26_E_T | inv_op_3 & _tlb_26_E_T_2 | inv_op_4
     & _tlb_26_E_T_5 | inv_op_5 & _tlb_26_E_T_8;
  wire  _tlb_27_E_T = ~tlb_27_G;
  wire  _tlb_27_E_T_2 = _tlb_27_E_T & asidMatch_27_1;
  wire  _tlb_27_E_T_5 = _tlb_27_E_T_2 & vaMatch_27_1;
  wire  _tlb_27_E_T_8 = (_tlb_27_E_T | asidMatch_27_1) & vaMatch_27_1;
  wire  _tlb_27_E_T_19 = inv_op_0 | inv_op_1 & tlb_27_G | inv_op_2 & _tlb_27_E_T | inv_op_3 & _tlb_27_E_T_2 | inv_op_4
     & _tlb_27_E_T_5 | inv_op_5 & _tlb_27_E_T_8;
  wire  _tlb_28_E_T = ~tlb_28_G;
  wire  _tlb_28_E_T_2 = _tlb_28_E_T & asidMatch_28_1;
  wire  _tlb_28_E_T_5 = _tlb_28_E_T_2 & vaMatch_28_1;
  wire  _tlb_28_E_T_8 = (_tlb_28_E_T | asidMatch_28_1) & vaMatch_28_1;
  wire  _tlb_28_E_T_19 = inv_op_0 | inv_op_1 & tlb_28_G | inv_op_2 & _tlb_28_E_T | inv_op_3 & _tlb_28_E_T_2 | inv_op_4
     & _tlb_28_E_T_5 | inv_op_5 & _tlb_28_E_T_8;
  wire  _tlb_29_E_T = ~tlb_29_G;
  wire  _tlb_29_E_T_2 = _tlb_29_E_T & asidMatch_29_1;
  wire  _tlb_29_E_T_5 = _tlb_29_E_T_2 & vaMatch_29_1;
  wire  _tlb_29_E_T_8 = (_tlb_29_E_T | asidMatch_29_1) & vaMatch_29_1;
  wire  _tlb_29_E_T_19 = inv_op_0 | inv_op_1 & tlb_29_G | inv_op_2 & _tlb_29_E_T | inv_op_3 & _tlb_29_E_T_2 | inv_op_4
     & _tlb_29_E_T_5 | inv_op_5 & _tlb_29_E_T_8;
  wire  _tlb_30_E_T = ~tlb_30_G;
  wire  _tlb_30_E_T_2 = _tlb_30_E_T & asidMatch_30_1;
  wire  _tlb_30_E_T_5 = _tlb_30_E_T_2 & vaMatch_30_1;
  wire  _tlb_30_E_T_8 = (_tlb_30_E_T | asidMatch_30_1) & vaMatch_30_1;
  wire  _tlb_30_E_T_19 = inv_op_0 | inv_op_1 & tlb_30_G | inv_op_2 & _tlb_30_E_T | inv_op_3 & _tlb_30_E_T_2 | inv_op_4
     & _tlb_30_E_T_5 | inv_op_5 & _tlb_30_E_T_8;
  wire  _tlb_31_E_T = ~tlb_31_G;
  wire  _tlb_31_E_T_2 = _tlb_31_E_T & asidMatch_31_1;
  wire  _tlb_31_E_T_5 = _tlb_31_E_T_2 & vaMatch_31_1;
  wire  _tlb_31_E_T_8 = (_tlb_31_E_T | asidMatch_31_1) & vaMatch_31_1;
  wire  _tlb_31_E_T_19 = inv_op_0 | inv_op_1 & tlb_31_G | inv_op_2 & _tlb_31_E_T | inv_op_3 & _tlb_31_E_T_2 | inv_op_4
     & _tlb_31_E_T_5 | inv_op_5 & _tlb_31_E_T_8;
  wire  _GEN_1745 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_0_E & ~_tlb_0_E_T_19 : tlb_0_E
    ;
  wire  _GEN_1746 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_1_E & ~_tlb_1_E_T_19 : tlb_1_E
    ;
  wire  _GEN_1747 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_2_E & ~_tlb_2_E_T_19 : tlb_2_E
    ;
  wire  _GEN_1748 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_3_E & ~_tlb_3_E_T_19 : tlb_3_E
    ;
  wire  _GEN_1749 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_4_E & ~_tlb_4_E_T_19 : tlb_4_E
    ;
  wire  _GEN_1750 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_5_E & ~_tlb_5_E_T_19 : tlb_5_E
    ;
  wire  _GEN_1751 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_6_E & ~_tlb_6_E_T_19 : tlb_6_E
    ;
  wire  _GEN_1752 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_7_E & ~_tlb_7_E_T_19 : tlb_7_E
    ;
  wire  _GEN_1753 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_8_E & ~_tlb_8_E_T_19 : tlb_8_E
    ;
  wire  _GEN_1754 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_9_E & ~_tlb_9_E_T_19 : tlb_9_E
    ;
  wire  _GEN_1755 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_10_E & ~_tlb_10_E_T_19 :
    tlb_10_E;
  wire  _GEN_1756 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_11_E & ~_tlb_11_E_T_19 :
    tlb_11_E;
  wire  _GEN_1757 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_12_E & ~_tlb_12_E_T_19 :
    tlb_12_E;
  wire  _GEN_1758 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_13_E & ~_tlb_13_E_T_19 :
    tlb_13_E;
  wire  _GEN_1759 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_14_E & ~_tlb_14_E_T_19 :
    tlb_14_E;
  wire  _GEN_1760 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_15_E & ~_tlb_15_E_T_19 :
    tlb_15_E;
  wire  _GEN_1761 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_16_E & ~_tlb_16_E_T_19 :
    tlb_16_E;
  wire  _GEN_1762 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_17_E & ~_tlb_17_E_T_19 :
    tlb_17_E;
  wire  _GEN_1763 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_18_E & ~_tlb_18_E_T_19 :
    tlb_18_E;
  wire  _GEN_1764 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_19_E & ~_tlb_19_E_T_19 :
    tlb_19_E;
  wire  _GEN_1765 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_20_E & ~_tlb_20_E_T_19 :
    tlb_20_E;
  wire  _GEN_1766 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_21_E & ~_tlb_21_E_T_19 :
    tlb_21_E;
  wire  _GEN_1767 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_22_E & ~_tlb_22_E_T_19 :
    tlb_22_E;
  wire  _GEN_1768 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_23_E & ~_tlb_23_E_T_19 :
    tlb_23_E;
  wire  _GEN_1769 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_24_E & ~_tlb_24_E_T_19 :
    tlb_24_E;
  wire  _GEN_1770 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_25_E & ~_tlb_25_E_T_19 :
    tlb_25_E;
  wire  _GEN_1771 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_26_E & ~_tlb_26_E_T_19 :
    tlb_26_E;
  wire  _GEN_1772 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_27_E & ~_tlb_27_E_T_19 :
    tlb_27_E;
  wire  _GEN_1773 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_28_E & ~_tlb_28_E_T_19 :
    tlb_28_E;
  wire  _GEN_1774 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_29_E & ~_tlb_29_E_T_19 :
    tlb_29_E;
  wire  _GEN_1775 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_30_E & ~_tlb_30_E_T_19 :
    tlb_30_E;
  wire  _GEN_1776 = inv_op_0 | inv_op_1 | inv_op_2 | inv_op_3 | inv_op_4 | inv_op_5 ? tlb_31_E & ~_tlb_31_E_T_19 :
    tlb_31_E;
  wire  _GEN_1778 = _T_1479 ? _GEN_1745 : tlb_0_E;
  wire  _GEN_1779 = _T_1479 ? _GEN_1746 : tlb_1_E;
  wire  _GEN_1780 = _T_1479 ? _GEN_1747 : tlb_2_E;
  wire  _GEN_1781 = _T_1479 ? _GEN_1748 : tlb_3_E;
  wire  _GEN_1782 = _T_1479 ? _GEN_1749 : tlb_4_E;
  wire  _GEN_1783 = _T_1479 ? _GEN_1750 : tlb_5_E;
  wire  _GEN_1784 = _T_1479 ? _GEN_1751 : tlb_6_E;
  wire  _GEN_1785 = _T_1479 ? _GEN_1752 : tlb_7_E;
  wire  _GEN_1786 = _T_1479 ? _GEN_1753 : tlb_8_E;
  wire  _GEN_1787 = _T_1479 ? _GEN_1754 : tlb_9_E;
  wire  _GEN_1788 = _T_1479 ? _GEN_1755 : tlb_10_E;
  wire  _GEN_1789 = _T_1479 ? _GEN_1756 : tlb_11_E;
  wire  _GEN_1790 = _T_1479 ? _GEN_1757 : tlb_12_E;
  wire  _GEN_1791 = _T_1479 ? _GEN_1758 : tlb_13_E;
  wire  _GEN_1792 = _T_1479 ? _GEN_1759 : tlb_14_E;
  wire  _GEN_1793 = _T_1479 ? _GEN_1760 : tlb_15_E;
  wire  _GEN_1794 = _T_1479 ? _GEN_1761 : tlb_16_E;
  wire  _GEN_1795 = _T_1479 ? _GEN_1762 : tlb_17_E;
  wire  _GEN_1796 = _T_1479 ? _GEN_1763 : tlb_18_E;
  wire  _GEN_1797 = _T_1479 ? _GEN_1764 : tlb_19_E;
  wire  _GEN_1798 = _T_1479 ? _GEN_1765 : tlb_20_E;
  wire  _GEN_1799 = _T_1479 ? _GEN_1766 : tlb_21_E;
  wire  _GEN_1800 = _T_1479 ? _GEN_1767 : tlb_22_E;
  wire  _GEN_1801 = _T_1479 ? _GEN_1768 : tlb_23_E;
  wire  _GEN_1802 = _T_1479 ? _GEN_1769 : tlb_24_E;
  wire  _GEN_1803 = _T_1479 ? _GEN_1770 : tlb_25_E;
  wire  _GEN_1804 = _T_1479 ? _GEN_1771 : tlb_26_E;
  wire  _GEN_1805 = _T_1479 ? _GEN_1772 : tlb_27_E;
  wire  _GEN_1806 = _T_1479 ? _GEN_1773 : tlb_28_E;
  wire  _GEN_1807 = _T_1479 ? _GEN_1774 : tlb_29_E;
  wire  _GEN_1808 = _T_1479 ? _GEN_1775 : tlb_30_E;
  wire  _GEN_1809 = _T_1479 ? _GEN_1776 : tlb_31_E;
  wire [18:0] _GEN_1811 = _T_1477 ? _GEN_1265 : tlb_0_VPPN;
  wire [18:0] _GEN_1812 = _T_1477 ? _GEN_1266 : tlb_1_VPPN;
  wire [18:0] _GEN_1813 = _T_1477 ? _GEN_1267 : tlb_2_VPPN;
  wire [18:0] _GEN_1814 = _T_1477 ? _GEN_1268 : tlb_3_VPPN;
  wire [18:0] _GEN_1815 = _T_1477 ? _GEN_1269 : tlb_4_VPPN;
  wire [18:0] _GEN_1816 = _T_1477 ? _GEN_1270 : tlb_5_VPPN;
  wire [18:0] _GEN_1817 = _T_1477 ? _GEN_1271 : tlb_6_VPPN;
  wire [18:0] _GEN_1818 = _T_1477 ? _GEN_1272 : tlb_7_VPPN;
  wire [18:0] _GEN_1819 = _T_1477 ? _GEN_1273 : tlb_8_VPPN;
  wire [18:0] _GEN_1820 = _T_1477 ? _GEN_1274 : tlb_9_VPPN;
  wire [18:0] _GEN_1821 = _T_1477 ? _GEN_1275 : tlb_10_VPPN;
  wire [18:0] _GEN_1822 = _T_1477 ? _GEN_1276 : tlb_11_VPPN;
  wire [18:0] _GEN_1823 = _T_1477 ? _GEN_1277 : tlb_12_VPPN;
  wire [18:0] _GEN_1824 = _T_1477 ? _GEN_1278 : tlb_13_VPPN;
  wire [18:0] _GEN_1825 = _T_1477 ? _GEN_1279 : tlb_14_VPPN;
  wire [18:0] _GEN_1826 = _T_1477 ? _GEN_1280 : tlb_15_VPPN;
  wire [18:0] _GEN_1827 = _T_1477 ? _GEN_1281 : tlb_16_VPPN;
  wire [18:0] _GEN_1828 = _T_1477 ? _GEN_1282 : tlb_17_VPPN;
  wire [18:0] _GEN_1829 = _T_1477 ? _GEN_1283 : tlb_18_VPPN;
  wire [18:0] _GEN_1830 = _T_1477 ? _GEN_1284 : tlb_19_VPPN;
  wire [18:0] _GEN_1831 = _T_1477 ? _GEN_1285 : tlb_20_VPPN;
  wire [18:0] _GEN_1832 = _T_1477 ? _GEN_1286 : tlb_21_VPPN;
  wire [18:0] _GEN_1833 = _T_1477 ? _GEN_1287 : tlb_22_VPPN;
  wire [18:0] _GEN_1834 = _T_1477 ? _GEN_1288 : tlb_23_VPPN;
  wire [18:0] _GEN_1835 = _T_1477 ? _GEN_1289 : tlb_24_VPPN;
  wire [18:0] _GEN_1836 = _T_1477 ? _GEN_1290 : tlb_25_VPPN;
  wire [18:0] _GEN_1837 = _T_1477 ? _GEN_1291 : tlb_26_VPPN;
  wire [18:0] _GEN_1838 = _T_1477 ? _GEN_1292 : tlb_27_VPPN;
  wire [18:0] _GEN_1839 = _T_1477 ? _GEN_1293 : tlb_28_VPPN;
  wire [18:0] _GEN_1840 = _T_1477 ? _GEN_1294 : tlb_29_VPPN;
  wire [18:0] _GEN_1841 = _T_1477 ? _GEN_1295 : tlb_30_VPPN;
  wire [18:0] _GEN_1842 = _T_1477 ? _GEN_1296 : tlb_31_VPPN;
  wire [5:0] _GEN_1843 = _T_1477 ? _GEN_1297 : tlb_0_PS;
  wire [5:0] _GEN_1844 = _T_1477 ? _GEN_1298 : tlb_1_PS;
  wire [5:0] _GEN_1845 = _T_1477 ? _GEN_1299 : tlb_2_PS;
  wire [5:0] _GEN_1846 = _T_1477 ? _GEN_1300 : tlb_3_PS;
  wire [5:0] _GEN_1847 = _T_1477 ? _GEN_1301 : tlb_4_PS;
  wire [5:0] _GEN_1848 = _T_1477 ? _GEN_1302 : tlb_5_PS;
  wire [5:0] _GEN_1849 = _T_1477 ? _GEN_1303 : tlb_6_PS;
  wire [5:0] _GEN_1850 = _T_1477 ? _GEN_1304 : tlb_7_PS;
  wire [5:0] _GEN_1851 = _T_1477 ? _GEN_1305 : tlb_8_PS;
  wire [5:0] _GEN_1852 = _T_1477 ? _GEN_1306 : tlb_9_PS;
  wire [5:0] _GEN_1853 = _T_1477 ? _GEN_1307 : tlb_10_PS;
  wire [5:0] _GEN_1854 = _T_1477 ? _GEN_1308 : tlb_11_PS;
  wire [5:0] _GEN_1855 = _T_1477 ? _GEN_1309 : tlb_12_PS;
  wire [5:0] _GEN_1856 = _T_1477 ? _GEN_1310 : tlb_13_PS;
  wire [5:0] _GEN_1857 = _T_1477 ? _GEN_1311 : tlb_14_PS;
  wire [5:0] _GEN_1858 = _T_1477 ? _GEN_1312 : tlb_15_PS;
  wire [5:0] _GEN_1859 = _T_1477 ? _GEN_1313 : tlb_16_PS;
  wire [5:0] _GEN_1860 = _T_1477 ? _GEN_1314 : tlb_17_PS;
  wire [5:0] _GEN_1861 = _T_1477 ? _GEN_1315 : tlb_18_PS;
  wire [5:0] _GEN_1862 = _T_1477 ? _GEN_1316 : tlb_19_PS;
  wire [5:0] _GEN_1863 = _T_1477 ? _GEN_1317 : tlb_20_PS;
  wire [5:0] _GEN_1864 = _T_1477 ? _GEN_1318 : tlb_21_PS;
  wire [5:0] _GEN_1865 = _T_1477 ? _GEN_1319 : tlb_22_PS;
  wire [5:0] _GEN_1866 = _T_1477 ? _GEN_1320 : tlb_23_PS;
  wire [5:0] _GEN_1867 = _T_1477 ? _GEN_1321 : tlb_24_PS;
  wire [5:0] _GEN_1868 = _T_1477 ? _GEN_1322 : tlb_25_PS;
  wire [5:0] _GEN_1869 = _T_1477 ? _GEN_1323 : tlb_26_PS;
  wire [5:0] _GEN_1870 = _T_1477 ? _GEN_1324 : tlb_27_PS;
  wire [5:0] _GEN_1871 = _T_1477 ? _GEN_1325 : tlb_28_PS;
  wire [5:0] _GEN_1872 = _T_1477 ? _GEN_1326 : tlb_29_PS;
  wire [5:0] _GEN_1873 = _T_1477 ? _GEN_1327 : tlb_30_PS;
  wire [5:0] _GEN_1874 = _T_1477 ? _GEN_1328 : tlb_31_PS;
  wire  _GEN_1875 = _T_1477 ? _GEN_1329 : tlb_0_G;
  wire  _GEN_1876 = _T_1477 ? _GEN_1330 : tlb_1_G;
  wire  _GEN_1877 = _T_1477 ? _GEN_1331 : tlb_2_G;
  wire  _GEN_1878 = _T_1477 ? _GEN_1332 : tlb_3_G;
  wire  _GEN_1879 = _T_1477 ? _GEN_1333 : tlb_4_G;
  wire  _GEN_1880 = _T_1477 ? _GEN_1334 : tlb_5_G;
  wire  _GEN_1881 = _T_1477 ? _GEN_1335 : tlb_6_G;
  wire  _GEN_1882 = _T_1477 ? _GEN_1336 : tlb_7_G;
  wire  _GEN_1883 = _T_1477 ? _GEN_1337 : tlb_8_G;
  wire  _GEN_1884 = _T_1477 ? _GEN_1338 : tlb_9_G;
  wire  _GEN_1885 = _T_1477 ? _GEN_1339 : tlb_10_G;
  wire  _GEN_1886 = _T_1477 ? _GEN_1340 : tlb_11_G;
  wire  _GEN_1887 = _T_1477 ? _GEN_1341 : tlb_12_G;
  wire  _GEN_1888 = _T_1477 ? _GEN_1342 : tlb_13_G;
  wire  _GEN_1889 = _T_1477 ? _GEN_1343 : tlb_14_G;
  wire  _GEN_1890 = _T_1477 ? _GEN_1344 : tlb_15_G;
  wire  _GEN_1891 = _T_1477 ? _GEN_1345 : tlb_16_G;
  wire  _GEN_1892 = _T_1477 ? _GEN_1346 : tlb_17_G;
  wire  _GEN_1893 = _T_1477 ? _GEN_1347 : tlb_18_G;
  wire  _GEN_1894 = _T_1477 ? _GEN_1348 : tlb_19_G;
  wire  _GEN_1895 = _T_1477 ? _GEN_1349 : tlb_20_G;
  wire  _GEN_1896 = _T_1477 ? _GEN_1350 : tlb_21_G;
  wire  _GEN_1897 = _T_1477 ? _GEN_1351 : tlb_22_G;
  wire  _GEN_1898 = _T_1477 ? _GEN_1352 : tlb_23_G;
  wire  _GEN_1899 = _T_1477 ? _GEN_1353 : tlb_24_G;
  wire  _GEN_1900 = _T_1477 ? _GEN_1354 : tlb_25_G;
  wire  _GEN_1901 = _T_1477 ? _GEN_1355 : tlb_26_G;
  wire  _GEN_1902 = _T_1477 ? _GEN_1356 : tlb_27_G;
  wire  _GEN_1903 = _T_1477 ? _GEN_1357 : tlb_28_G;
  wire  _GEN_1904 = _T_1477 ? _GEN_1358 : tlb_29_G;
  wire  _GEN_1905 = _T_1477 ? _GEN_1359 : tlb_30_G;
  wire  _GEN_1906 = _T_1477 ? _GEN_1360 : tlb_31_G;
  wire [9:0] _GEN_1907 = _T_1477 ? _GEN_1361 : tlb_0_ASID;
  wire [9:0] _GEN_1908 = _T_1477 ? _GEN_1362 : tlb_1_ASID;
  wire [9:0] _GEN_1909 = _T_1477 ? _GEN_1363 : tlb_2_ASID;
  wire [9:0] _GEN_1910 = _T_1477 ? _GEN_1364 : tlb_3_ASID;
  wire [9:0] _GEN_1911 = _T_1477 ? _GEN_1365 : tlb_4_ASID;
  wire [9:0] _GEN_1912 = _T_1477 ? _GEN_1366 : tlb_5_ASID;
  wire [9:0] _GEN_1913 = _T_1477 ? _GEN_1367 : tlb_6_ASID;
  wire [9:0] _GEN_1914 = _T_1477 ? _GEN_1368 : tlb_7_ASID;
  wire [9:0] _GEN_1915 = _T_1477 ? _GEN_1369 : tlb_8_ASID;
  wire [9:0] _GEN_1916 = _T_1477 ? _GEN_1370 : tlb_9_ASID;
  wire [9:0] _GEN_1917 = _T_1477 ? _GEN_1371 : tlb_10_ASID;
  wire [9:0] _GEN_1918 = _T_1477 ? _GEN_1372 : tlb_11_ASID;
  wire [9:0] _GEN_1919 = _T_1477 ? _GEN_1373 : tlb_12_ASID;
  wire [9:0] _GEN_1920 = _T_1477 ? _GEN_1374 : tlb_13_ASID;
  wire [9:0] _GEN_1921 = _T_1477 ? _GEN_1375 : tlb_14_ASID;
  wire [9:0] _GEN_1922 = _T_1477 ? _GEN_1376 : tlb_15_ASID;
  wire [9:0] _GEN_1923 = _T_1477 ? _GEN_1377 : tlb_16_ASID;
  wire [9:0] _GEN_1924 = _T_1477 ? _GEN_1378 : tlb_17_ASID;
  wire [9:0] _GEN_1925 = _T_1477 ? _GEN_1379 : tlb_18_ASID;
  wire [9:0] _GEN_1926 = _T_1477 ? _GEN_1380 : tlb_19_ASID;
  wire [9:0] _GEN_1927 = _T_1477 ? _GEN_1381 : tlb_20_ASID;
  wire [9:0] _GEN_1928 = _T_1477 ? _GEN_1382 : tlb_21_ASID;
  wire [9:0] _GEN_1929 = _T_1477 ? _GEN_1383 : tlb_22_ASID;
  wire [9:0] _GEN_1930 = _T_1477 ? _GEN_1384 : tlb_23_ASID;
  wire [9:0] _GEN_1931 = _T_1477 ? _GEN_1385 : tlb_24_ASID;
  wire [9:0] _GEN_1932 = _T_1477 ? _GEN_1386 : tlb_25_ASID;
  wire [9:0] _GEN_1933 = _T_1477 ? _GEN_1387 : tlb_26_ASID;
  wire [9:0] _GEN_1934 = _T_1477 ? _GEN_1388 : tlb_27_ASID;
  wire [9:0] _GEN_1935 = _T_1477 ? _GEN_1389 : tlb_28_ASID;
  wire [9:0] _GEN_1936 = _T_1477 ? _GEN_1390 : tlb_29_ASID;
  wire [9:0] _GEN_1937 = _T_1477 ? _GEN_1391 : tlb_30_ASID;
  wire [9:0] _GEN_1938 = _T_1477 ? _GEN_1392 : tlb_31_ASID;
  wire  _GEN_1939 = _T_1477 ? _GEN_1393 : _GEN_1778;
  wire  _GEN_1940 = _T_1477 ? _GEN_1394 : _GEN_1779;
  wire  _GEN_1941 = _T_1477 ? _GEN_1395 : _GEN_1780;
  wire  _GEN_1942 = _T_1477 ? _GEN_1396 : _GEN_1781;
  wire  _GEN_1943 = _T_1477 ? _GEN_1397 : _GEN_1782;
  wire  _GEN_1944 = _T_1477 ? _GEN_1398 : _GEN_1783;
  wire  _GEN_1945 = _T_1477 ? _GEN_1399 : _GEN_1784;
  wire  _GEN_1946 = _T_1477 ? _GEN_1400 : _GEN_1785;
  wire  _GEN_1947 = _T_1477 ? _GEN_1401 : _GEN_1786;
  wire  _GEN_1948 = _T_1477 ? _GEN_1402 : _GEN_1787;
  wire  _GEN_1949 = _T_1477 ? _GEN_1403 : _GEN_1788;
  wire  _GEN_1950 = _T_1477 ? _GEN_1404 : _GEN_1789;
  wire  _GEN_1951 = _T_1477 ? _GEN_1405 : _GEN_1790;
  wire  _GEN_1952 = _T_1477 ? _GEN_1406 : _GEN_1791;
  wire  _GEN_1953 = _T_1477 ? _GEN_1407 : _GEN_1792;
  wire  _GEN_1954 = _T_1477 ? _GEN_1408 : _GEN_1793;
  wire  _GEN_1955 = _T_1477 ? _GEN_1409 : _GEN_1794;
  wire  _GEN_1956 = _T_1477 ? _GEN_1410 : _GEN_1795;
  wire  _GEN_1957 = _T_1477 ? _GEN_1411 : _GEN_1796;
  wire  _GEN_1958 = _T_1477 ? _GEN_1412 : _GEN_1797;
  wire  _GEN_1959 = _T_1477 ? _GEN_1413 : _GEN_1798;
  wire  _GEN_1960 = _T_1477 ? _GEN_1414 : _GEN_1799;
  wire  _GEN_1961 = _T_1477 ? _GEN_1415 : _GEN_1800;
  wire  _GEN_1962 = _T_1477 ? _GEN_1416 : _GEN_1801;
  wire  _GEN_1963 = _T_1477 ? _GEN_1417 : _GEN_1802;
  wire  _GEN_1964 = _T_1477 ? _GEN_1418 : _GEN_1803;
  wire  _GEN_1965 = _T_1477 ? _GEN_1419 : _GEN_1804;
  wire  _GEN_1966 = _T_1477 ? _GEN_1420 : _GEN_1805;
  wire  _GEN_1967 = _T_1477 ? _GEN_1421 : _GEN_1806;
  wire  _GEN_1968 = _T_1477 ? _GEN_1422 : _GEN_1807;
  wire  _GEN_1969 = _T_1477 ? _GEN_1423 : _GEN_1808;
  wire  _GEN_1970 = _T_1477 ? _GEN_1424 : _GEN_1809;
  wire [19:0] _GEN_1971 = _T_1477 ? _GEN_1425 : tlb_0_P0_PPN;
  wire [19:0] _GEN_1972 = _T_1477 ? _GEN_1426 : tlb_1_P0_PPN;
  wire [19:0] _GEN_1973 = _T_1477 ? _GEN_1427 : tlb_2_P0_PPN;
  wire [19:0] _GEN_1974 = _T_1477 ? _GEN_1428 : tlb_3_P0_PPN;
  wire [19:0] _GEN_1975 = _T_1477 ? _GEN_1429 : tlb_4_P0_PPN;
  wire [19:0] _GEN_1976 = _T_1477 ? _GEN_1430 : tlb_5_P0_PPN;
  wire [19:0] _GEN_1977 = _T_1477 ? _GEN_1431 : tlb_6_P0_PPN;
  wire [19:0] _GEN_1978 = _T_1477 ? _GEN_1432 : tlb_7_P0_PPN;
  wire [19:0] _GEN_1979 = _T_1477 ? _GEN_1433 : tlb_8_P0_PPN;
  wire [19:0] _GEN_1980 = _T_1477 ? _GEN_1434 : tlb_9_P0_PPN;
  wire [19:0] _GEN_1981 = _T_1477 ? _GEN_1435 : tlb_10_P0_PPN;
  wire [19:0] _GEN_1982 = _T_1477 ? _GEN_1436 : tlb_11_P0_PPN;
  wire [19:0] _GEN_1983 = _T_1477 ? _GEN_1437 : tlb_12_P0_PPN;
  wire [19:0] _GEN_1984 = _T_1477 ? _GEN_1438 : tlb_13_P0_PPN;
  wire [19:0] _GEN_1985 = _T_1477 ? _GEN_1439 : tlb_14_P0_PPN;
  wire [19:0] _GEN_1986 = _T_1477 ? _GEN_1440 : tlb_15_P0_PPN;
  wire [19:0] _GEN_1987 = _T_1477 ? _GEN_1441 : tlb_16_P0_PPN;
  wire [19:0] _GEN_1988 = _T_1477 ? _GEN_1442 : tlb_17_P0_PPN;
  wire [19:0] _GEN_1989 = _T_1477 ? _GEN_1443 : tlb_18_P0_PPN;
  wire [19:0] _GEN_1990 = _T_1477 ? _GEN_1444 : tlb_19_P0_PPN;
  wire [19:0] _GEN_1991 = _T_1477 ? _GEN_1445 : tlb_20_P0_PPN;
  wire [19:0] _GEN_1992 = _T_1477 ? _GEN_1446 : tlb_21_P0_PPN;
  wire [19:0] _GEN_1993 = _T_1477 ? _GEN_1447 : tlb_22_P0_PPN;
  wire [19:0] _GEN_1994 = _T_1477 ? _GEN_1448 : tlb_23_P0_PPN;
  wire [19:0] _GEN_1995 = _T_1477 ? _GEN_1449 : tlb_24_P0_PPN;
  wire [19:0] _GEN_1996 = _T_1477 ? _GEN_1450 : tlb_25_P0_PPN;
  wire [19:0] _GEN_1997 = _T_1477 ? _GEN_1451 : tlb_26_P0_PPN;
  wire [19:0] _GEN_1998 = _T_1477 ? _GEN_1452 : tlb_27_P0_PPN;
  wire [19:0] _GEN_1999 = _T_1477 ? _GEN_1453 : tlb_28_P0_PPN;
  wire [19:0] _GEN_2000 = _T_1477 ? _GEN_1454 : tlb_29_P0_PPN;
  wire [19:0] _GEN_2001 = _T_1477 ? _GEN_1455 : tlb_30_P0_PPN;
  wire [19:0] _GEN_2002 = _T_1477 ? _GEN_1456 : tlb_31_P0_PPN;
  wire [1:0] _GEN_2003 = _T_1477 ? _GEN_1457 : tlb_0_P0_PLV;
  wire [1:0] _GEN_2004 = _T_1477 ? _GEN_1458 : tlb_1_P0_PLV;
  wire [1:0] _GEN_2005 = _T_1477 ? _GEN_1459 : tlb_2_P0_PLV;
  wire [1:0] _GEN_2006 = _T_1477 ? _GEN_1460 : tlb_3_P0_PLV;
  wire [1:0] _GEN_2007 = _T_1477 ? _GEN_1461 : tlb_4_P0_PLV;
  wire [1:0] _GEN_2008 = _T_1477 ? _GEN_1462 : tlb_5_P0_PLV;
  wire [1:0] _GEN_2009 = _T_1477 ? _GEN_1463 : tlb_6_P0_PLV;
  wire [1:0] _GEN_2010 = _T_1477 ? _GEN_1464 : tlb_7_P0_PLV;
  wire [1:0] _GEN_2011 = _T_1477 ? _GEN_1465 : tlb_8_P0_PLV;
  wire [1:0] _GEN_2012 = _T_1477 ? _GEN_1466 : tlb_9_P0_PLV;
  wire [1:0] _GEN_2013 = _T_1477 ? _GEN_1467 : tlb_10_P0_PLV;
  wire [1:0] _GEN_2014 = _T_1477 ? _GEN_1468 : tlb_11_P0_PLV;
  wire [1:0] _GEN_2015 = _T_1477 ? _GEN_1469 : tlb_12_P0_PLV;
  wire [1:0] _GEN_2016 = _T_1477 ? _GEN_1470 : tlb_13_P0_PLV;
  wire [1:0] _GEN_2017 = _T_1477 ? _GEN_1471 : tlb_14_P0_PLV;
  wire [1:0] _GEN_2018 = _T_1477 ? _GEN_1472 : tlb_15_P0_PLV;
  wire [1:0] _GEN_2019 = _T_1477 ? _GEN_1473 : tlb_16_P0_PLV;
  wire [1:0] _GEN_2020 = _T_1477 ? _GEN_1474 : tlb_17_P0_PLV;
  wire [1:0] _GEN_2021 = _T_1477 ? _GEN_1475 : tlb_18_P0_PLV;
  wire [1:0] _GEN_2022 = _T_1477 ? _GEN_1476 : tlb_19_P0_PLV;
  wire [1:0] _GEN_2023 = _T_1477 ? _GEN_1477 : tlb_20_P0_PLV;
  wire [1:0] _GEN_2024 = _T_1477 ? _GEN_1478 : tlb_21_P0_PLV;
  wire [1:0] _GEN_2025 = _T_1477 ? _GEN_1479 : tlb_22_P0_PLV;
  wire [1:0] _GEN_2026 = _T_1477 ? _GEN_1480 : tlb_23_P0_PLV;
  wire [1:0] _GEN_2027 = _T_1477 ? _GEN_1481 : tlb_24_P0_PLV;
  wire [1:0] _GEN_2028 = _T_1477 ? _GEN_1482 : tlb_25_P0_PLV;
  wire [1:0] _GEN_2029 = _T_1477 ? _GEN_1483 : tlb_26_P0_PLV;
  wire [1:0] _GEN_2030 = _T_1477 ? _GEN_1484 : tlb_27_P0_PLV;
  wire [1:0] _GEN_2031 = _T_1477 ? _GEN_1485 : tlb_28_P0_PLV;
  wire [1:0] _GEN_2032 = _T_1477 ? _GEN_1486 : tlb_29_P0_PLV;
  wire [1:0] _GEN_2033 = _T_1477 ? _GEN_1487 : tlb_30_P0_PLV;
  wire [1:0] _GEN_2034 = _T_1477 ? _GEN_1488 : tlb_31_P0_PLV;
  wire [1:0] _GEN_2035 = _T_1477 ? _GEN_1489 : tlb_0_P0_MAT;
  wire [1:0] _GEN_2036 = _T_1477 ? _GEN_1490 : tlb_1_P0_MAT;
  wire [1:0] _GEN_2037 = _T_1477 ? _GEN_1491 : tlb_2_P0_MAT;
  wire [1:0] _GEN_2038 = _T_1477 ? _GEN_1492 : tlb_3_P0_MAT;
  wire [1:0] _GEN_2039 = _T_1477 ? _GEN_1493 : tlb_4_P0_MAT;
  wire [1:0] _GEN_2040 = _T_1477 ? _GEN_1494 : tlb_5_P0_MAT;
  wire [1:0] _GEN_2041 = _T_1477 ? _GEN_1495 : tlb_6_P0_MAT;
  wire [1:0] _GEN_2042 = _T_1477 ? _GEN_1496 : tlb_7_P0_MAT;
  wire [1:0] _GEN_2043 = _T_1477 ? _GEN_1497 : tlb_8_P0_MAT;
  wire [1:0] _GEN_2044 = _T_1477 ? _GEN_1498 : tlb_9_P0_MAT;
  wire [1:0] _GEN_2045 = _T_1477 ? _GEN_1499 : tlb_10_P0_MAT;
  wire [1:0] _GEN_2046 = _T_1477 ? _GEN_1500 : tlb_11_P0_MAT;
  wire [1:0] _GEN_2047 = _T_1477 ? _GEN_1501 : tlb_12_P0_MAT;
  wire [1:0] _GEN_2048 = _T_1477 ? _GEN_1502 : tlb_13_P0_MAT;
  wire [1:0] _GEN_2049 = _T_1477 ? _GEN_1503 : tlb_14_P0_MAT;
  wire [1:0] _GEN_2050 = _T_1477 ? _GEN_1504 : tlb_15_P0_MAT;
  wire [1:0] _GEN_2051 = _T_1477 ? _GEN_1505 : tlb_16_P0_MAT;
  wire [1:0] _GEN_2052 = _T_1477 ? _GEN_1506 : tlb_17_P0_MAT;
  wire [1:0] _GEN_2053 = _T_1477 ? _GEN_1507 : tlb_18_P0_MAT;
  wire [1:0] _GEN_2054 = _T_1477 ? _GEN_1508 : tlb_19_P0_MAT;
  wire [1:0] _GEN_2055 = _T_1477 ? _GEN_1509 : tlb_20_P0_MAT;
  wire [1:0] _GEN_2056 = _T_1477 ? _GEN_1510 : tlb_21_P0_MAT;
  wire [1:0] _GEN_2057 = _T_1477 ? _GEN_1511 : tlb_22_P0_MAT;
  wire [1:0] _GEN_2058 = _T_1477 ? _GEN_1512 : tlb_23_P0_MAT;
  wire [1:0] _GEN_2059 = _T_1477 ? _GEN_1513 : tlb_24_P0_MAT;
  wire [1:0] _GEN_2060 = _T_1477 ? _GEN_1514 : tlb_25_P0_MAT;
  wire [1:0] _GEN_2061 = _T_1477 ? _GEN_1515 : tlb_26_P0_MAT;
  wire [1:0] _GEN_2062 = _T_1477 ? _GEN_1516 : tlb_27_P0_MAT;
  wire [1:0] _GEN_2063 = _T_1477 ? _GEN_1517 : tlb_28_P0_MAT;
  wire [1:0] _GEN_2064 = _T_1477 ? _GEN_1518 : tlb_29_P0_MAT;
  wire [1:0] _GEN_2065 = _T_1477 ? _GEN_1519 : tlb_30_P0_MAT;
  wire [1:0] _GEN_2066 = _T_1477 ? _GEN_1520 : tlb_31_P0_MAT;
  wire  _GEN_2067 = _T_1477 ? _GEN_1521 : tlb_0_P0_D;
  wire  _GEN_2068 = _T_1477 ? _GEN_1522 : tlb_1_P0_D;
  wire  _GEN_2069 = _T_1477 ? _GEN_1523 : tlb_2_P0_D;
  wire  _GEN_2070 = _T_1477 ? _GEN_1524 : tlb_3_P0_D;
  wire  _GEN_2071 = _T_1477 ? _GEN_1525 : tlb_4_P0_D;
  wire  _GEN_2072 = _T_1477 ? _GEN_1526 : tlb_5_P0_D;
  wire  _GEN_2073 = _T_1477 ? _GEN_1527 : tlb_6_P0_D;
  wire  _GEN_2074 = _T_1477 ? _GEN_1528 : tlb_7_P0_D;
  wire  _GEN_2075 = _T_1477 ? _GEN_1529 : tlb_8_P0_D;
  wire  _GEN_2076 = _T_1477 ? _GEN_1530 : tlb_9_P0_D;
  wire  _GEN_2077 = _T_1477 ? _GEN_1531 : tlb_10_P0_D;
  wire  _GEN_2078 = _T_1477 ? _GEN_1532 : tlb_11_P0_D;
  wire  _GEN_2079 = _T_1477 ? _GEN_1533 : tlb_12_P0_D;
  wire  _GEN_2080 = _T_1477 ? _GEN_1534 : tlb_13_P0_D;
  wire  _GEN_2081 = _T_1477 ? _GEN_1535 : tlb_14_P0_D;
  wire  _GEN_2082 = _T_1477 ? _GEN_1536 : tlb_15_P0_D;
  wire  _GEN_2083 = _T_1477 ? _GEN_1537 : tlb_16_P0_D;
  wire  _GEN_2084 = _T_1477 ? _GEN_1538 : tlb_17_P0_D;
  wire  _GEN_2085 = _T_1477 ? _GEN_1539 : tlb_18_P0_D;
  wire  _GEN_2086 = _T_1477 ? _GEN_1540 : tlb_19_P0_D;
  wire  _GEN_2087 = _T_1477 ? _GEN_1541 : tlb_20_P0_D;
  wire  _GEN_2088 = _T_1477 ? _GEN_1542 : tlb_21_P0_D;
  wire  _GEN_2089 = _T_1477 ? _GEN_1543 : tlb_22_P0_D;
  wire  _GEN_2090 = _T_1477 ? _GEN_1544 : tlb_23_P0_D;
  wire  _GEN_2091 = _T_1477 ? _GEN_1545 : tlb_24_P0_D;
  wire  _GEN_2092 = _T_1477 ? _GEN_1546 : tlb_25_P0_D;
  wire  _GEN_2093 = _T_1477 ? _GEN_1547 : tlb_26_P0_D;
  wire  _GEN_2094 = _T_1477 ? _GEN_1548 : tlb_27_P0_D;
  wire  _GEN_2095 = _T_1477 ? _GEN_1549 : tlb_28_P0_D;
  wire  _GEN_2096 = _T_1477 ? _GEN_1550 : tlb_29_P0_D;
  wire  _GEN_2097 = _T_1477 ? _GEN_1551 : tlb_30_P0_D;
  wire  _GEN_2098 = _T_1477 ? _GEN_1552 : tlb_31_P0_D;
  wire  _GEN_2099 = _T_1477 ? _GEN_1553 : tlb_0_P0_V;
  wire  _GEN_2100 = _T_1477 ? _GEN_1554 : tlb_1_P0_V;
  wire  _GEN_2101 = _T_1477 ? _GEN_1555 : tlb_2_P0_V;
  wire  _GEN_2102 = _T_1477 ? _GEN_1556 : tlb_3_P0_V;
  wire  _GEN_2103 = _T_1477 ? _GEN_1557 : tlb_4_P0_V;
  wire  _GEN_2104 = _T_1477 ? _GEN_1558 : tlb_5_P0_V;
  wire  _GEN_2105 = _T_1477 ? _GEN_1559 : tlb_6_P0_V;
  wire  _GEN_2106 = _T_1477 ? _GEN_1560 : tlb_7_P0_V;
  wire  _GEN_2107 = _T_1477 ? _GEN_1561 : tlb_8_P0_V;
  wire  _GEN_2108 = _T_1477 ? _GEN_1562 : tlb_9_P0_V;
  wire  _GEN_2109 = _T_1477 ? _GEN_1563 : tlb_10_P0_V;
  wire  _GEN_2110 = _T_1477 ? _GEN_1564 : tlb_11_P0_V;
  wire  _GEN_2111 = _T_1477 ? _GEN_1565 : tlb_12_P0_V;
  wire  _GEN_2112 = _T_1477 ? _GEN_1566 : tlb_13_P0_V;
  wire  _GEN_2113 = _T_1477 ? _GEN_1567 : tlb_14_P0_V;
  wire  _GEN_2114 = _T_1477 ? _GEN_1568 : tlb_15_P0_V;
  wire  _GEN_2115 = _T_1477 ? _GEN_1569 : tlb_16_P0_V;
  wire  _GEN_2116 = _T_1477 ? _GEN_1570 : tlb_17_P0_V;
  wire  _GEN_2117 = _T_1477 ? _GEN_1571 : tlb_18_P0_V;
  wire  _GEN_2118 = _T_1477 ? _GEN_1572 : tlb_19_P0_V;
  wire  _GEN_2119 = _T_1477 ? _GEN_1573 : tlb_20_P0_V;
  wire  _GEN_2120 = _T_1477 ? _GEN_1574 : tlb_21_P0_V;
  wire  _GEN_2121 = _T_1477 ? _GEN_1575 : tlb_22_P0_V;
  wire  _GEN_2122 = _T_1477 ? _GEN_1576 : tlb_23_P0_V;
  wire  _GEN_2123 = _T_1477 ? _GEN_1577 : tlb_24_P0_V;
  wire  _GEN_2124 = _T_1477 ? _GEN_1578 : tlb_25_P0_V;
  wire  _GEN_2125 = _T_1477 ? _GEN_1579 : tlb_26_P0_V;
  wire  _GEN_2126 = _T_1477 ? _GEN_1580 : tlb_27_P0_V;
  wire  _GEN_2127 = _T_1477 ? _GEN_1581 : tlb_28_P0_V;
  wire  _GEN_2128 = _T_1477 ? _GEN_1582 : tlb_29_P0_V;
  wire  _GEN_2129 = _T_1477 ? _GEN_1583 : tlb_30_P0_V;
  wire  _GEN_2130 = _T_1477 ? _GEN_1584 : tlb_31_P0_V;
  wire [19:0] _GEN_2131 = _T_1477 ? _GEN_1585 : tlb_0_P1_PPN;
  wire [19:0] _GEN_2132 = _T_1477 ? _GEN_1586 : tlb_1_P1_PPN;
  wire [19:0] _GEN_2133 = _T_1477 ? _GEN_1587 : tlb_2_P1_PPN;
  wire [19:0] _GEN_2134 = _T_1477 ? _GEN_1588 : tlb_3_P1_PPN;
  wire [19:0] _GEN_2135 = _T_1477 ? _GEN_1589 : tlb_4_P1_PPN;
  wire [19:0] _GEN_2136 = _T_1477 ? _GEN_1590 : tlb_5_P1_PPN;
  wire [19:0] _GEN_2137 = _T_1477 ? _GEN_1591 : tlb_6_P1_PPN;
  wire [19:0] _GEN_2138 = _T_1477 ? _GEN_1592 : tlb_7_P1_PPN;
  wire [19:0] _GEN_2139 = _T_1477 ? _GEN_1593 : tlb_8_P1_PPN;
  wire [19:0] _GEN_2140 = _T_1477 ? _GEN_1594 : tlb_9_P1_PPN;
  wire [19:0] _GEN_2141 = _T_1477 ? _GEN_1595 : tlb_10_P1_PPN;
  wire [19:0] _GEN_2142 = _T_1477 ? _GEN_1596 : tlb_11_P1_PPN;
  wire [19:0] _GEN_2143 = _T_1477 ? _GEN_1597 : tlb_12_P1_PPN;
  wire [19:0] _GEN_2144 = _T_1477 ? _GEN_1598 : tlb_13_P1_PPN;
  wire [19:0] _GEN_2145 = _T_1477 ? _GEN_1599 : tlb_14_P1_PPN;
  wire [19:0] _GEN_2146 = _T_1477 ? _GEN_1600 : tlb_15_P1_PPN;
  wire [19:0] _GEN_2147 = _T_1477 ? _GEN_1601 : tlb_16_P1_PPN;
  wire [19:0] _GEN_2148 = _T_1477 ? _GEN_1602 : tlb_17_P1_PPN;
  wire [19:0] _GEN_2149 = _T_1477 ? _GEN_1603 : tlb_18_P1_PPN;
  wire [19:0] _GEN_2150 = _T_1477 ? _GEN_1604 : tlb_19_P1_PPN;
  wire [19:0] _GEN_2151 = _T_1477 ? _GEN_1605 : tlb_20_P1_PPN;
  wire [19:0] _GEN_2152 = _T_1477 ? _GEN_1606 : tlb_21_P1_PPN;
  wire [19:0] _GEN_2153 = _T_1477 ? _GEN_1607 : tlb_22_P1_PPN;
  wire [19:0] _GEN_2154 = _T_1477 ? _GEN_1608 : tlb_23_P1_PPN;
  wire [19:0] _GEN_2155 = _T_1477 ? _GEN_1609 : tlb_24_P1_PPN;
  wire [19:0] _GEN_2156 = _T_1477 ? _GEN_1610 : tlb_25_P1_PPN;
  wire [19:0] _GEN_2157 = _T_1477 ? _GEN_1611 : tlb_26_P1_PPN;
  wire [19:0] _GEN_2158 = _T_1477 ? _GEN_1612 : tlb_27_P1_PPN;
  wire [19:0] _GEN_2159 = _T_1477 ? _GEN_1613 : tlb_28_P1_PPN;
  wire [19:0] _GEN_2160 = _T_1477 ? _GEN_1614 : tlb_29_P1_PPN;
  wire [19:0] _GEN_2161 = _T_1477 ? _GEN_1615 : tlb_30_P1_PPN;
  wire [19:0] _GEN_2162 = _T_1477 ? _GEN_1616 : tlb_31_P1_PPN;
  wire [1:0] _GEN_2163 = _T_1477 ? _GEN_1617 : tlb_0_P1_PLV;
  wire [1:0] _GEN_2164 = _T_1477 ? _GEN_1618 : tlb_1_P1_PLV;
  wire [1:0] _GEN_2165 = _T_1477 ? _GEN_1619 : tlb_2_P1_PLV;
  wire [1:0] _GEN_2166 = _T_1477 ? _GEN_1620 : tlb_3_P1_PLV;
  wire [1:0] _GEN_2167 = _T_1477 ? _GEN_1621 : tlb_4_P1_PLV;
  wire [1:0] _GEN_2168 = _T_1477 ? _GEN_1622 : tlb_5_P1_PLV;
  wire [1:0] _GEN_2169 = _T_1477 ? _GEN_1623 : tlb_6_P1_PLV;
  wire [1:0] _GEN_2170 = _T_1477 ? _GEN_1624 : tlb_7_P1_PLV;
  wire [1:0] _GEN_2171 = _T_1477 ? _GEN_1625 : tlb_8_P1_PLV;
  wire [1:0] _GEN_2172 = _T_1477 ? _GEN_1626 : tlb_9_P1_PLV;
  wire [1:0] _GEN_2173 = _T_1477 ? _GEN_1627 : tlb_10_P1_PLV;
  wire [1:0] _GEN_2174 = _T_1477 ? _GEN_1628 : tlb_11_P1_PLV;
  wire [1:0] _GEN_2175 = _T_1477 ? _GEN_1629 : tlb_12_P1_PLV;
  wire [1:0] _GEN_2176 = _T_1477 ? _GEN_1630 : tlb_13_P1_PLV;
  wire [1:0] _GEN_2177 = _T_1477 ? _GEN_1631 : tlb_14_P1_PLV;
  wire [1:0] _GEN_2178 = _T_1477 ? _GEN_1632 : tlb_15_P1_PLV;
  wire [1:0] _GEN_2179 = _T_1477 ? _GEN_1633 : tlb_16_P1_PLV;
  wire [1:0] _GEN_2180 = _T_1477 ? _GEN_1634 : tlb_17_P1_PLV;
  wire [1:0] _GEN_2181 = _T_1477 ? _GEN_1635 : tlb_18_P1_PLV;
  wire [1:0] _GEN_2182 = _T_1477 ? _GEN_1636 : tlb_19_P1_PLV;
  wire [1:0] _GEN_2183 = _T_1477 ? _GEN_1637 : tlb_20_P1_PLV;
  wire [1:0] _GEN_2184 = _T_1477 ? _GEN_1638 : tlb_21_P1_PLV;
  wire [1:0] _GEN_2185 = _T_1477 ? _GEN_1639 : tlb_22_P1_PLV;
  wire [1:0] _GEN_2186 = _T_1477 ? _GEN_1640 : tlb_23_P1_PLV;
  wire [1:0] _GEN_2187 = _T_1477 ? _GEN_1641 : tlb_24_P1_PLV;
  wire [1:0] _GEN_2188 = _T_1477 ? _GEN_1642 : tlb_25_P1_PLV;
  wire [1:0] _GEN_2189 = _T_1477 ? _GEN_1643 : tlb_26_P1_PLV;
  wire [1:0] _GEN_2190 = _T_1477 ? _GEN_1644 : tlb_27_P1_PLV;
  wire [1:0] _GEN_2191 = _T_1477 ? _GEN_1645 : tlb_28_P1_PLV;
  wire [1:0] _GEN_2192 = _T_1477 ? _GEN_1646 : tlb_29_P1_PLV;
  wire [1:0] _GEN_2193 = _T_1477 ? _GEN_1647 : tlb_30_P1_PLV;
  wire [1:0] _GEN_2194 = _T_1477 ? _GEN_1648 : tlb_31_P1_PLV;
  wire [1:0] _GEN_2195 = _T_1477 ? _GEN_1649 : tlb_0_P1_MAT;
  wire [1:0] _GEN_2196 = _T_1477 ? _GEN_1650 : tlb_1_P1_MAT;
  wire [1:0] _GEN_2197 = _T_1477 ? _GEN_1651 : tlb_2_P1_MAT;
  wire [1:0] _GEN_2198 = _T_1477 ? _GEN_1652 : tlb_3_P1_MAT;
  wire [1:0] _GEN_2199 = _T_1477 ? _GEN_1653 : tlb_4_P1_MAT;
  wire [1:0] _GEN_2200 = _T_1477 ? _GEN_1654 : tlb_5_P1_MAT;
  wire [1:0] _GEN_2201 = _T_1477 ? _GEN_1655 : tlb_6_P1_MAT;
  wire [1:0] _GEN_2202 = _T_1477 ? _GEN_1656 : tlb_7_P1_MAT;
  wire [1:0] _GEN_2203 = _T_1477 ? _GEN_1657 : tlb_8_P1_MAT;
  wire [1:0] _GEN_2204 = _T_1477 ? _GEN_1658 : tlb_9_P1_MAT;
  wire [1:0] _GEN_2205 = _T_1477 ? _GEN_1659 : tlb_10_P1_MAT;
  wire [1:0] _GEN_2206 = _T_1477 ? _GEN_1660 : tlb_11_P1_MAT;
  wire [1:0] _GEN_2207 = _T_1477 ? _GEN_1661 : tlb_12_P1_MAT;
  wire [1:0] _GEN_2208 = _T_1477 ? _GEN_1662 : tlb_13_P1_MAT;
  wire [1:0] _GEN_2209 = _T_1477 ? _GEN_1663 : tlb_14_P1_MAT;
  wire [1:0] _GEN_2210 = _T_1477 ? _GEN_1664 : tlb_15_P1_MAT;
  wire [1:0] _GEN_2211 = _T_1477 ? _GEN_1665 : tlb_16_P1_MAT;
  wire [1:0] _GEN_2212 = _T_1477 ? _GEN_1666 : tlb_17_P1_MAT;
  wire [1:0] _GEN_2213 = _T_1477 ? _GEN_1667 : tlb_18_P1_MAT;
  wire [1:0] _GEN_2214 = _T_1477 ? _GEN_1668 : tlb_19_P1_MAT;
  wire [1:0] _GEN_2215 = _T_1477 ? _GEN_1669 : tlb_20_P1_MAT;
  wire [1:0] _GEN_2216 = _T_1477 ? _GEN_1670 : tlb_21_P1_MAT;
  wire [1:0] _GEN_2217 = _T_1477 ? _GEN_1671 : tlb_22_P1_MAT;
  wire [1:0] _GEN_2218 = _T_1477 ? _GEN_1672 : tlb_23_P1_MAT;
  wire [1:0] _GEN_2219 = _T_1477 ? _GEN_1673 : tlb_24_P1_MAT;
  wire [1:0] _GEN_2220 = _T_1477 ? _GEN_1674 : tlb_25_P1_MAT;
  wire [1:0] _GEN_2221 = _T_1477 ? _GEN_1675 : tlb_26_P1_MAT;
  wire [1:0] _GEN_2222 = _T_1477 ? _GEN_1676 : tlb_27_P1_MAT;
  wire [1:0] _GEN_2223 = _T_1477 ? _GEN_1677 : tlb_28_P1_MAT;
  wire [1:0] _GEN_2224 = _T_1477 ? _GEN_1678 : tlb_29_P1_MAT;
  wire [1:0] _GEN_2225 = _T_1477 ? _GEN_1679 : tlb_30_P1_MAT;
  wire [1:0] _GEN_2226 = _T_1477 ? _GEN_1680 : tlb_31_P1_MAT;
  wire  _GEN_2227 = _T_1477 ? _GEN_1681 : tlb_0_P1_D;
  wire  _GEN_2228 = _T_1477 ? _GEN_1682 : tlb_1_P1_D;
  wire  _GEN_2229 = _T_1477 ? _GEN_1683 : tlb_2_P1_D;
  wire  _GEN_2230 = _T_1477 ? _GEN_1684 : tlb_3_P1_D;
  wire  _GEN_2231 = _T_1477 ? _GEN_1685 : tlb_4_P1_D;
  wire  _GEN_2232 = _T_1477 ? _GEN_1686 : tlb_5_P1_D;
  wire  _GEN_2233 = _T_1477 ? _GEN_1687 : tlb_6_P1_D;
  wire  _GEN_2234 = _T_1477 ? _GEN_1688 : tlb_7_P1_D;
  wire  _GEN_2235 = _T_1477 ? _GEN_1689 : tlb_8_P1_D;
  wire  _GEN_2236 = _T_1477 ? _GEN_1690 : tlb_9_P1_D;
  wire  _GEN_2237 = _T_1477 ? _GEN_1691 : tlb_10_P1_D;
  wire  _GEN_2238 = _T_1477 ? _GEN_1692 : tlb_11_P1_D;
  wire  _GEN_2239 = _T_1477 ? _GEN_1693 : tlb_12_P1_D;
  wire  _GEN_2240 = _T_1477 ? _GEN_1694 : tlb_13_P1_D;
  wire  _GEN_2241 = _T_1477 ? _GEN_1695 : tlb_14_P1_D;
  wire  _GEN_2242 = _T_1477 ? _GEN_1696 : tlb_15_P1_D;
  wire  _GEN_2243 = _T_1477 ? _GEN_1697 : tlb_16_P1_D;
  wire  _GEN_2244 = _T_1477 ? _GEN_1698 : tlb_17_P1_D;
  wire  _GEN_2245 = _T_1477 ? _GEN_1699 : tlb_18_P1_D;
  wire  _GEN_2246 = _T_1477 ? _GEN_1700 : tlb_19_P1_D;
  wire  _GEN_2247 = _T_1477 ? _GEN_1701 : tlb_20_P1_D;
  wire  _GEN_2248 = _T_1477 ? _GEN_1702 : tlb_21_P1_D;
  wire  _GEN_2249 = _T_1477 ? _GEN_1703 : tlb_22_P1_D;
  wire  _GEN_2250 = _T_1477 ? _GEN_1704 : tlb_23_P1_D;
  wire  _GEN_2251 = _T_1477 ? _GEN_1705 : tlb_24_P1_D;
  wire  _GEN_2252 = _T_1477 ? _GEN_1706 : tlb_25_P1_D;
  wire  _GEN_2253 = _T_1477 ? _GEN_1707 : tlb_26_P1_D;
  wire  _GEN_2254 = _T_1477 ? _GEN_1708 : tlb_27_P1_D;
  wire  _GEN_2255 = _T_1477 ? _GEN_1709 : tlb_28_P1_D;
  wire  _GEN_2256 = _T_1477 ? _GEN_1710 : tlb_29_P1_D;
  wire  _GEN_2257 = _T_1477 ? _GEN_1711 : tlb_30_P1_D;
  wire  _GEN_2258 = _T_1477 ? _GEN_1712 : tlb_31_P1_D;
  wire  _GEN_2259 = _T_1477 ? _GEN_1713 : tlb_0_P1_V;
  wire  _GEN_2260 = _T_1477 ? _GEN_1714 : tlb_1_P1_V;
  wire  _GEN_2261 = _T_1477 ? _GEN_1715 : tlb_2_P1_V;
  wire  _GEN_2262 = _T_1477 ? _GEN_1716 : tlb_3_P1_V;
  wire  _GEN_2263 = _T_1477 ? _GEN_1717 : tlb_4_P1_V;
  wire  _GEN_2264 = _T_1477 ? _GEN_1718 : tlb_5_P1_V;
  wire  _GEN_2265 = _T_1477 ? _GEN_1719 : tlb_6_P1_V;
  wire  _GEN_2266 = _T_1477 ? _GEN_1720 : tlb_7_P1_V;
  wire  _GEN_2267 = _T_1477 ? _GEN_1721 : tlb_8_P1_V;
  wire  _GEN_2268 = _T_1477 ? _GEN_1722 : tlb_9_P1_V;
  wire  _GEN_2269 = _T_1477 ? _GEN_1723 : tlb_10_P1_V;
  wire  _GEN_2270 = _T_1477 ? _GEN_1724 : tlb_11_P1_V;
  wire  _GEN_2271 = _T_1477 ? _GEN_1725 : tlb_12_P1_V;
  wire  _GEN_2272 = _T_1477 ? _GEN_1726 : tlb_13_P1_V;
  wire  _GEN_2273 = _T_1477 ? _GEN_1727 : tlb_14_P1_V;
  wire  _GEN_2274 = _T_1477 ? _GEN_1728 : tlb_15_P1_V;
  wire  _GEN_2275 = _T_1477 ? _GEN_1729 : tlb_16_P1_V;
  wire  _GEN_2276 = _T_1477 ? _GEN_1730 : tlb_17_P1_V;
  wire  _GEN_2277 = _T_1477 ? _GEN_1731 : tlb_18_P1_V;
  wire  _GEN_2278 = _T_1477 ? _GEN_1732 : tlb_19_P1_V;
  wire  _GEN_2279 = _T_1477 ? _GEN_1733 : tlb_20_P1_V;
  wire  _GEN_2280 = _T_1477 ? _GEN_1734 : tlb_21_P1_V;
  wire  _GEN_2281 = _T_1477 ? _GEN_1735 : tlb_22_P1_V;
  wire  _GEN_2282 = _T_1477 ? _GEN_1736 : tlb_23_P1_V;
  wire  _GEN_2283 = _T_1477 ? _GEN_1737 : tlb_24_P1_V;
  wire  _GEN_2284 = _T_1477 ? _GEN_1738 : tlb_25_P1_V;
  wire  _GEN_2285 = _T_1477 ? _GEN_1739 : tlb_26_P1_V;
  wire  _GEN_2286 = _T_1477 ? _GEN_1740 : tlb_27_P1_V;
  wire  _GEN_2287 = _T_1477 ? _GEN_1741 : tlb_28_P1_V;
  wire  _GEN_2288 = _T_1477 ? _GEN_1742 : tlb_29_P1_V;
  wire  _GEN_2289 = _T_1477 ? _GEN_1743 : tlb_30_P1_V;
  wire  _GEN_2290 = _T_1477 ? _GEN_1744 : tlb_31_P1_V;
  wire  _wbIdx_T_1 = c0_1 == 2'h1;
  wire  _wbIdx_T_2 = c0_1 == 2'h2;
  wire  _wbIdx_T_3 = c0_1 == 2'h3;
  wire [4:0] _wbIdx_T_5 = _wbIdx_T_1 ? 5'h1 : 5'h0;
  wire [4:0] _wbIdx_T_6 = _wbIdx_T_2 ? d : 5'h0;
  wire [4:0] _wbIdx_T_7 = _wbIdx_T_3 ? j : 5'h0;
  wire [4:0] _wbIdx_T_9 = _wbIdx_T_5 | _wbIdx_T_6;
  wire [4:0] wbIdx = _wbIdx_T_9 | _wbIdx_T_7;
  wire  _wbData_T = c0_0 == 3'h0;
  wire  _wbData_T_1 = c0_0 == 3'h1;
  wire  _wbData_T_2 = c0_0 == 3'h2;
  wire  _wbData_T_3 = c0_0 == 3'h3;
  wire  _wbData_T_4 = c0_0 == 3'h4;
  wire  _wbData_T_5 = c0_0 == 3'h5;
  wire  _wbData_T_7 = c0_0 == 3'h6;
  wire  _wbData_T_9 = c0_0 == 3'h7;
  wire [31:0] _wbData_T_10 = _wbData_T ? aluOut : 32'h0;
  wire [31:0] _wbData_T_11 = _wbData_T_1 ? extendData : 32'h0;
  wire [31:0] _wbData_T_12 = _wbData_T_2 ? PC4 : 32'h0;
  wire [31:0] _wbData_T_13 = _wbData_T_3 ? csrRD : 32'h0;
  wire [31:0] _wbData_T_14 = _wbData_T_4 ? csrs_21_TID : 32'h0;
  wire [31:0] _wbData_T_15 = _wbData_T_5 ? timer[63:32] : 32'h0;
  wire [31:0] _wbData_T_16 = _wbData_T_7 ? timer[31:0] : 32'h0;
  wire  _wbData_T_17 = _wbData_T_9 & csrs_25_ROLLB;
  wire [31:0] _wbData_T_18 = _wbData_T_10 | _wbData_T_11;
  wire [31:0] _wbData_T_19 = _wbData_T_18 | _wbData_T_12;
  wire [31:0] _wbData_T_20 = _wbData_T_19 | _wbData_T_13;
  wire [31:0] _wbData_T_21 = _wbData_T_20 | _wbData_T_14;
  wire [31:0] _wbData_T_22 = _wbData_T_21 | _wbData_T_15;
  wire [31:0] _wbData_T_23 = _wbData_T_22 | _wbData_T_16;
  wire [31:0] _GEN_4333 = {{31'd0}, _wbData_T_17};
  wire  _T_1486 = mem_OK & |wbIdx;
  wire  _T_1487 = ~dStall;
  wire  _GEN_4273 = _tlb_E_T | _GEN_234;
  wire  _GEN_4274 = _tlb_E_T ? 1'h0 : _GEN_233;
  wire [1:0] _GEN_4275 = ID_OK & c0_8 ? csrs_1_PPLV : _GEN_231;
  wire  _GEN_4276 = ID_OK & c0_8 ? csrs_1_PIE : _GEN_232;
  wire  _GEN_4279 = ID_OK & c0_8 ? _GEN_4273 : _GEN_234;
  wire  _GEN_4280 = ID_OK & c0_8 ? _GEN_4274 : _GEN_233;
  wire  _GEN_4281 = ID_OK & c0_9 | idle;
  wire  _T_1495 = _T_1319 & _T_1487;
  wire [3:0] _estat_Ecode_T_1 = ADEF ? 4'h8 : 4'h0;
  wire [1:0] _estat_Ecode_T_2 = PIF ? 2'h3 : 2'h0;
  wire [3:0] _estat_Ecode_T_3 = INE ? 4'hd : 4'h0;
  wire [3:0] _estat_Ecode_T_5 = SYS ? 4'hb : 4'h0;
  wire [3:0] _estat_Ecode_T_6 = BRK ? 4'hc : 4'h0;
  wire [3:0] _estat_Ecode_T_7 = ALE ? 4'h9 : 4'h0;
  wire [3:0] _estat_Ecode_T_8 = ADEM ? 4'h8 : 4'h0;
  wire [1:0] _estat_Ecode_T_10 = PIS ? 2'h2 : 2'h0;
  wire [2:0] _estat_Ecode_T_11 = PME ? 3'h4 : 3'h0;
  wire [2:0] _estat_Ecode_T_12 = PPI ? 3'h7 : 3'h0;
  wire [5:0] _estat_Ecode_T_15 = TLBR ? 6'h3f : 6'h0;
  wire [3:0] _GEN_4334 = {{2'd0}, _estat_Ecode_T_2};
  wire [3:0] _estat_Ecode_T_17 = _estat_Ecode_T_1 | _GEN_4334;
  wire [3:0] _estat_Ecode_T_18 = _estat_Ecode_T_17 | _estat_Ecode_T_3;
  wire [3:0] _estat_Ecode_T_20 = _estat_Ecode_T_18 | _estat_Ecode_T_5;
  wire [3:0] _estat_Ecode_T_21 = _estat_Ecode_T_20 | _estat_Ecode_T_6;
  wire [3:0] _estat_Ecode_T_22 = _estat_Ecode_T_21 | _estat_Ecode_T_7;
  wire [3:0] _estat_Ecode_T_23 = _estat_Ecode_T_22 | _estat_Ecode_T_8;
  wire [3:0] _GEN_4335 = {{3'd0}, PIL};
  wire [3:0] _estat_Ecode_T_24 = _estat_Ecode_T_23 | _GEN_4335;
  wire [3:0] _GEN_4336 = {{2'd0}, _estat_Ecode_T_10};
  wire [3:0] _estat_Ecode_T_25 = _estat_Ecode_T_24 | _GEN_4336;
  wire [3:0] _GEN_4337 = {{1'd0}, _estat_Ecode_T_11};
  wire [3:0] _estat_Ecode_T_26 = _estat_Ecode_T_25 | _GEN_4337;
  wire [3:0] _GEN_4338 = {{1'd0}, _estat_Ecode_T_12};
  wire [3:0] _estat_Ecode_T_27 = _estat_Ecode_T_26 | _GEN_4338;
  wire [4:0] _estat_Ecode_T_29 = {{1'd0}, _estat_Ecode_T_27};
  wire [5:0] _GEN_4339 = {{1'd0}, _estat_Ecode_T_29};
  wire [5:0] _estat_Ecode_T_30 = _GEN_4339 | _estat_Ecode_T_15;
  wire  _GEN_4290 = TLBR | _GEN_4280;
  wire  _GEN_4300 = _T_1319 & _T_1487 ? _GEN_4290 : _GEN_4280;
  wire  _take_T = rj != rkd;
  wire  _take_T_1 = rj == rkd;
  wire [31:0] _take_T_2 = j == 5'h0 ? 32'h0 : GR_rj_MPORT_data;
  wire [31:0] _take_T_3 = kd == 5'h0 ? 32'h0 : GR_rkd_MPORT_data;
  wire  _take_T_4 = $signed(_take_T_2) >= $signed(_take_T_3);
  wire  _take_T_5 = rj >= rkd;
  wire  _take_T_8 = $signed(_take_T_2) < $signed(_take_T_3);
  wire  _take_T_9 = rj < rkd;
  wire  _GEN_4304 = 3'h2 == brType ? _take_T_1 : 3'h1 == brType & _take_T;
  wire  _GEN_4305 = 3'h3 == brType ? _take_T_4 : _GEN_4304;
  wire  _GEN_4306 = 3'h4 == brType ? _take_T_5 : _GEN_4305;
  wire  _GEN_4307 = 3'h5 == brType ? _take_T_8 : _GEN_4306;
  wire  _GEN_4308 = 3'h6 == brType ? _take_T_9 : _GEN_4307;
  wire [31:0] _PC_T_2 = 3'h7 == brType | _GEN_4308 ? aluOut : PC4;
  wire [31:0] _GEN_4310 = _T_27 & ~(c0_9 & ID_OK) ? _PC_T_2 : PC;
  wire [31:0] _GEN_4311 = c0_8 ? csrs_5_PC : _GEN_4310;
  assign GR_rj_MPORT_addr = inst[9:5];
  assign GR_rj_MPORT_data = GR[GR_rj_MPORT_addr];
  assign GR_rkd_MPORT_addr = _kd_T_5 ? d : k;
  assign GR_rkd_MPORT_data = GR[GR_rkd_MPORT_addr];
  assign GR_MPORT_data = _wbData_T_23 | _GEN_4333;
  assign GR_MPORT_addr = _wbIdx_T_9 | _wbIdx_T_7;
  assign GR_MPORT_mask = 1'h1;
  assign GR_MPORT_en = _T_1486 & _T_1487;
  assign io_inst_req_valid = reset ? 1'h0 : ~iStallReg & ~dStallReg & IF_OK;
  assign io_inst_req_bits_addr = crmd_DA ? PC : pa;
  assign io_data_req_valid = reset ? 1'h0 : _io_inst_req_valid_T_1 & mem_OK & _EXVA_T & ~preldNop & ~(c0_11 & d[2:0] != 3'h1
    );
  assign io_data_req_bits_wen = _io_data_req_bits_wen_T_4[3:0];
  assign io_data_req_bits_addr = c0_11 & d[4:3] == 2'h2 | ~c0_11 & crmd_PG ? pa_1 : aluOut;
  assign io_data_req_bits_wdata = _io_data_req_bits_wdata_T_2[31:0];
  assign io_data_req_bits_cacop = _T_38 ? 1'h0 : _T_1254;
  assign io_data_req_bits_preld = _T_38 ? 1'h0 : _T_1318;
  assign io_debug_pc = PC;
  assign io_debug_wen = mem_OK & |wbIdx & ~dStall ? 4'hf : 4'h0;
  assign io_debug_wnum = _wbIdx_T_9 | _wbIdx_T_7;
  assign io_debug_wdata = _wbData_T_23 | _GEN_4333;
  always @(posedge clock) begin
    if(GR_MPORT_en & GR_MPORT_mask) begin
      GR[GR_MPORT_addr] <= GR_MPORT_data;
    end
    if (reset) begin
      idle <= 1'h0;
    end else if (_T_1319 & _T_1487) begin
      if (excp) begin
        idle <= 1'h0;
      end else begin
        idle <= _GEN_4281;
      end
    end else begin
      idle <= _GEN_4281;
    end
    if (reset) begin
      PC <= 32'h1c000000;
    end else if (_T_1495) begin
      if (TLBR) begin
        PC <= _csrRD_T_44;
      end else if (excp) begin
        PC <= _csrRD_T_11;
      end else begin
        PC <= _GEN_4311;
      end
    end
    if (reset) begin
      timer <= 64'h0;
    end else begin
      timer <= _timer_T_1;
    end
    if (reset) begin
      iStallReg <= 1'h0;
    end else begin
      iStallReg <= iStall;
    end
    if (reset) begin
      dStallReg <= 1'h0;
    end else begin
      dStallReg <= dStall;
    end
    if (reset) begin
      crmd_DATM <= 2'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T) begin
        crmd_DATM <= _crmd_T_4[8:7];
      end
    end
    if (reset) begin
      crmd_DATF <= 2'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T) begin
        crmd_DATF <= _crmd_T_4[6:5];
      end
    end
    if (reset) begin
      crmd_PG <= 1'h0;
    end else if (_T_1319 & _T_1487) begin
      if (TLBR) begin
        crmd_PG <= 1'h0;
      end else begin
        crmd_PG <= _GEN_4279;
      end
    end else begin
      crmd_PG <= _GEN_4279;
    end
    crmd_DA <= reset | _GEN_4300;
    if (reset) begin
      crmd_IE <= 1'h0;
    end else if (_T_1319 & _T_1487) begin
      if (excp) begin
        crmd_IE <= 1'h0;
      end else begin
        crmd_IE <= _GEN_4276;
      end
    end else begin
      crmd_IE <= _GEN_4276;
    end
    if (reset) begin
      crmd_PLV <= 2'h0;
    end else if (_T_1319 & _T_1487) begin
      if (excp) begin
        crmd_PLV <= 2'h0;
      end else begin
        crmd_PLV <= _GEN_4275;
      end
    end else begin
      crmd_PLV <= _GEN_4275;
    end
    if (reset) begin
      csrs_1_PIE <= 1'h0;
    end else if (_T_1319 & _T_1487) begin
      if (excp) begin
        csrs_1_PIE <= crmd_IE;
      end else begin
        csrs_1_PIE <= _GEN_238;
      end
    end else begin
      csrs_1_PIE <= _GEN_238;
    end
    if (reset) begin
      csrs_1_PPLV <= 2'h0;
    end else if (_T_1319 & _T_1487) begin
      if (excp) begin
        csrs_1_PPLV <= crmd_PLV;
      end else begin
        csrs_1_PPLV <= _GEN_237;
      end
    end else begin
      csrs_1_PPLV <= _GEN_237;
    end
    if (reset) begin
      csrs_2_FPE <= 1'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_4) begin
        csrs_2_FPE <= _euen_T_3[0];
      end
    end
    if (reset) begin
      csrs_3_LIE <= 13'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_5) begin
        csrs_3_LIE <= _ectl_T_3[12:0];
      end
    end
    if (reset) begin
      csrs_4_EsubCode <= 9'h0;
    end else if (_T_1319 & _T_1487) begin
      if (excp) begin
        csrs_4_EsubCode <= {{8'd0}, ADEM};
      end
    end
    if (reset) begin
      csrs_4_Ecode <= 6'h0;
    end else if (_T_1319 & _T_1487) begin
      if (excp) begin
        csrs_4_Ecode <= _estat_Ecode_T_30;
      end
    end
    if (reset) begin
      csrs_4_IS_0 <= 1'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_6) begin
        if (csrMask[0]) begin
          csrs_4_IS_0 <= rkd[0];
        end
      end
    end
    if (reset) begin
      csrs_4_IS_1 <= 1'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_6) begin
        if (csrMask[0]) begin
          csrs_4_IS_1 <= rkd[1];
        end
      end
    end
    if (reset) begin
      csrs_4_IS_2 <= 1'h0;
    end else begin
      csrs_4_IS_2 <= io_interrupt[0];
    end
    if (reset) begin
      csrs_4_IS_3 <= 1'h0;
    end else begin
      csrs_4_IS_3 <= io_interrupt[1];
    end
    if (reset) begin
      csrs_4_IS_4 <= 1'h0;
    end else begin
      csrs_4_IS_4 <= io_interrupt[2];
    end
    if (reset) begin
      csrs_4_IS_5 <= 1'h0;
    end else begin
      csrs_4_IS_5 <= io_interrupt[3];
    end
    if (reset) begin
      csrs_4_IS_6 <= 1'h0;
    end else begin
      csrs_4_IS_6 <= io_interrupt[4];
    end
    if (reset) begin
      csrs_4_IS_7 <= 1'h0;
    end else begin
      csrs_4_IS_7 <= io_interrupt[5];
    end
    if (reset) begin
      csrs_4_IS_8 <= 1'h0;
    end else begin
      csrs_4_IS_8 <= io_interrupt[6];
    end
    if (reset) begin
      csrs_4_IS_9 <= 1'h0;
    end else begin
      csrs_4_IS_9 <= io_interrupt[7];
    end
    if (reset) begin
      csrs_4_IS_11 <= 1'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_40) begin
        if (rkd[0] & csrMask[0]) begin
          csrs_4_IS_11 <= 1'h0;
        end else begin
          csrs_4_IS_11 <= _GEN_6;
        end
      end else begin
        csrs_4_IS_11 <= _GEN_6;
      end
    end else begin
      csrs_4_IS_11 <= _GEN_6;
    end
    if (reset) begin
      csrs_4_IS_12 <= 1'h0;
    end else begin
      csrs_4_IS_12 <= io_ipi;
    end
    if (reset) begin
      csrs_5_PC <= 32'h0;
    end else if (_T_1319 & _T_1487) begin
      if (excp) begin
        csrs_5_PC <= PC;
      end else begin
        csrs_5_PC <= _GEN_243;
      end
    end else begin
      csrs_5_PC <= _GEN_243;
    end
    if (reset) begin
      badv_VAddr <= 32'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_9) begin
        badv_VAddr <= _badv_T_3;
      end else begin
        badv_VAddr <= _GEN_167;
      end
    end else begin
      badv_VAddr <= _GEN_167;
    end
    if (reset) begin
      csrs_7_VA <= 26'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_10) begin
        csrs_7_VA <= _eentry_VA_T_3;
      end
    end
    if (reset) begin
      csrs_8_NE <= 1'h0;
    end else if (ID_OK) begin
      if (_T_1443) begin
        if (_miss_T_62) begin
          csrs_8_NE <= 1'h0;
        end else begin
          csrs_8_NE <= 1'h1;
        end
      end else if (_T_1475) begin
        csrs_8_NE <= ~_GEN_321;
      end else begin
        csrs_8_NE <= _GEN_246;
      end
    end else begin
      csrs_8_NE <= _GEN_246;
    end
    if (reset) begin
      csrs_8_PS <= 6'h0;
    end else if (ID_OK) begin
      if (_T_1443) begin
        csrs_8_PS <= _GEN_247;
      end else if (_T_1475) begin
        csrs_8_PS <= _GEN_770;
      end else begin
        csrs_8_PS <= _GEN_247;
      end
    end else begin
      csrs_8_PS <= _GEN_247;
    end
    if (reset) begin
      csrs_8_Index <= 5'h0;
    end else if (ID_OK) begin
      if (_T_1443) begin
        if (_miss_T_62) begin
          csrs_8_Index <= _tlbidx_Index_T_66;
        end else begin
          csrs_8_Index <= _GEN_248;
        end
      end else begin
        csrs_8_Index <= _GEN_248;
      end
    end else begin
      csrs_8_Index <= _GEN_248;
    end
    if (reset) begin
      csrs_9_VPPN <= 19'h0;
    end else if (ID_OK) begin
      if (_T_1443) begin
        csrs_9_VPPN <= _GEN_249;
      end else if (_T_1475) begin
        csrs_9_VPPN <= _GEN_771;
      end else begin
        csrs_9_VPPN <= _GEN_249;
      end
    end else begin
      csrs_9_VPPN <= _GEN_249;
    end
    if (reset) begin
      csrs_10_PPN <= 24'h0;
    end else if (ID_OK) begin
      if (_T_1443) begin
        csrs_10_PPN <= _GEN_255;
      end else if (_T_1475) begin
        csrs_10_PPN <= _GEN_772;
      end else begin
        csrs_10_PPN <= _GEN_255;
      end
    end else begin
      csrs_10_PPN <= _GEN_255;
    end
    if (reset) begin
      csrs_10_G <= 1'h0;
    end else if (ID_OK) begin
      if (_T_1443) begin
        csrs_10_G <= _GEN_254;
      end else if (_T_1475) begin
        csrs_10_G <= _GEN_773;
      end else begin
        csrs_10_G <= _GEN_254;
      end
    end else begin
      csrs_10_G <= _GEN_254;
    end
    if (reset) begin
      csrs_10_MAT <= 2'h0;
    end else if (ID_OK) begin
      if (_T_1443) begin
        csrs_10_MAT <= _GEN_253;
      end else if (_T_1475) begin
        csrs_10_MAT <= _GEN_774;
      end else begin
        csrs_10_MAT <= _GEN_253;
      end
    end else begin
      csrs_10_MAT <= _GEN_253;
    end
    if (reset) begin
      csrs_10_PLV <= 2'h0;
    end else if (ID_OK) begin
      if (_T_1443) begin
        csrs_10_PLV <= _GEN_252;
      end else if (_T_1475) begin
        csrs_10_PLV <= _GEN_775;
      end else begin
        csrs_10_PLV <= _GEN_252;
      end
    end else begin
      csrs_10_PLV <= _GEN_252;
    end
    if (reset) begin
      csrs_10_D <= 1'h0;
    end else if (ID_OK) begin
      if (_T_1443) begin
        csrs_10_D <= _GEN_251;
      end else if (_T_1475) begin
        csrs_10_D <= _GEN_776;
      end else begin
        csrs_10_D <= _GEN_251;
      end
    end else begin
      csrs_10_D <= _GEN_251;
    end
    if (reset) begin
      csrs_10_V <= 1'h0;
    end else if (ID_OK) begin
      if (_T_1443) begin
        csrs_10_V <= _GEN_250;
      end else if (_T_1475) begin
        csrs_10_V <= _GEN_777;
      end else begin
        csrs_10_V <= _GEN_250;
      end
    end else begin
      csrs_10_V <= _GEN_250;
    end
    if (reset) begin
      csrs_11_PPN <= 24'h0;
    end else if (ID_OK) begin
      if (_T_1443) begin
        csrs_11_PPN <= _GEN_261;
      end else if (_T_1475) begin
        csrs_11_PPN <= _GEN_778;
      end else begin
        csrs_11_PPN <= _GEN_261;
      end
    end else begin
      csrs_11_PPN <= _GEN_261;
    end
    if (reset) begin
      csrs_11_G <= 1'h0;
    end else if (ID_OK) begin
      if (_T_1443) begin
        csrs_11_G <= _GEN_260;
      end else if (_T_1475) begin
        csrs_11_G <= _GEN_779;
      end else begin
        csrs_11_G <= _GEN_260;
      end
    end else begin
      csrs_11_G <= _GEN_260;
    end
    if (reset) begin
      csrs_11_MAT <= 2'h0;
    end else if (ID_OK) begin
      if (_T_1443) begin
        csrs_11_MAT <= _GEN_259;
      end else if (_T_1475) begin
        csrs_11_MAT <= _GEN_780;
      end else begin
        csrs_11_MAT <= _GEN_259;
      end
    end else begin
      csrs_11_MAT <= _GEN_259;
    end
    if (reset) begin
      csrs_11_PLV <= 2'h0;
    end else if (ID_OK) begin
      if (_T_1443) begin
        csrs_11_PLV <= _GEN_258;
      end else if (_T_1475) begin
        csrs_11_PLV <= _GEN_781;
      end else begin
        csrs_11_PLV <= _GEN_258;
      end
    end else begin
      csrs_11_PLV <= _GEN_258;
    end
    if (reset) begin
      csrs_11_D <= 1'h0;
    end else if (ID_OK) begin
      if (_T_1443) begin
        csrs_11_D <= _GEN_257;
      end else if (_T_1475) begin
        csrs_11_D <= _GEN_782;
      end else begin
        csrs_11_D <= _GEN_257;
      end
    end else begin
      csrs_11_D <= _GEN_257;
    end
    if (reset) begin
      csrs_11_V <= 1'h0;
    end else if (ID_OK) begin
      if (_T_1443) begin
        csrs_11_V <= _GEN_256;
      end else if (_T_1475) begin
        csrs_11_V <= _GEN_783;
      end else begin
        csrs_11_V <= _GEN_256;
      end
    end else begin
      csrs_11_V <= _GEN_256;
    end
    if (reset) begin
      asid_ASID <= 10'h0;
    end else if (ID_OK) begin
      if (_T_1443) begin
        asid_ASID <= _GEN_262;
      end else if (_T_1475) begin
        asid_ASID <= _GEN_784;
      end else begin
        asid_ASID <= _GEN_262;
      end
    end else begin
      asid_ASID <= _GEN_262;
    end
    if (reset) begin
      csrs_13_Base <= 20'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_22) begin
        csrs_13_Base <= _pgdl_Base_T_3;
      end
    end
    if (reset) begin
      csrs_14_Base <= 20'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_24) begin
        csrs_14_Base <= _pgdh_Base_T_3;
      end
    end
    if (reset) begin
      csrs_17_Data <= 32'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_32) begin
        csrs_17_Data <= _save0_T_3;
      end
    end
    if (reset) begin
      csrs_18_Data <= 32'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_33) begin
        csrs_18_Data <= _save1_T_3;
      end
    end
    if (reset) begin
      csrs_19_Data <= 32'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_34) begin
        csrs_19_Data <= _save2_T_3;
      end
    end
    if (reset) begin
      csrs_20_Data <= 32'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_35) begin
        csrs_20_Data <= _save3_T_3;
      end
    end
    if (reset) begin
      csrs_21_TID <= 32'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_36) begin
        csrs_21_TID <= _tid_T_3;
      end
    end
    if (reset) begin
      csrs_22_InitVal <= 30'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_37) begin
        csrs_22_InitVal <= _tcfg_T_4[31:2];
      end
    end
    if (reset) begin
      csrs_22_Periodic <= 1'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_37) begin
        csrs_22_Periodic <= _tcfg_T_4[1];
      end
    end
    if (reset) begin
      csrs_22_En <= 1'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_37) begin
        csrs_22_En <= _tcfg_T_4[0];
      end else begin
        csrs_22_En <= _GEN_7;
      end
    end else begin
      csrs_22_En <= _GEN_7;
    end
    if (reset) begin
      csrs_23_TimeVal <= 32'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_37) begin
        csrs_23_TimeVal <= _tval_TimeVal_T_6;
      end else begin
        csrs_23_TimeVal <= _GEN_5;
      end
    end else begin
      csrs_23_TimeVal <= _GEN_5;
    end
    if (reset) begin
      csrs_25_KLO <= 1'h0;
    end else if (ID_OK & c0_8) begin
      csrs_25_KLO <= 1'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_41) begin
        csrs_25_KLO <= _GEN_216;
      end
    end
    if (reset) begin
      csrs_25_ROLLB <= 1'h0;
    end else if (ID_OK & c0_8) begin
      if (~csrs_25_KLO) begin
        csrs_25_ROLLB <= 1'h0;
      end else begin
        csrs_25_ROLLB <= _GEN_276;
      end
    end else begin
      csrs_25_ROLLB <= _GEN_276;
    end
    if (reset) begin
      csrs_26_PA <= 26'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_43) begin
        csrs_26_PA <= _tlbrentry_PA_T_3;
      end
    end
    if (reset) begin
      csrs_27_VSEG <= 3'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_45) begin
        csrs_27_VSEG <= _dmw0_VSEG_T_3;
      end
    end
    if (reset) begin
      csrs_27_PSEG <= 3'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_45) begin
        csrs_27_PSEG <= _dmw0_PSEG_T_3;
      end
    end
    if (reset) begin
      csrs_27_MAT <= 2'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_45) begin
        csrs_27_MAT <= _dmw0_MAT_T_3;
      end
    end
    if (reset) begin
      csrs_27_PLV3 <= 1'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_45) begin
        csrs_27_PLV3 <= rkd[3] & csrMask[3] | csrs_27_PLV3 & ~csrMask[3];
      end
    end
    if (reset) begin
      csrs_27_PLV0 <= 1'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_45) begin
        csrs_27_PLV0 <= _T_1412 | csrs_27_PLV0 & ~csrMask[0];
      end
    end
    if (reset) begin
      csrs_28_VSEG <= 3'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_47) begin
        csrs_28_VSEG <= _dmw1_VSEG_T_3;
      end
    end
    if (reset) begin
      csrs_28_PSEG <= 3'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_47) begin
        csrs_28_PSEG <= _dmw1_PSEG_T_3;
      end
    end
    if (reset) begin
      csrs_28_MAT <= 2'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_47) begin
        csrs_28_MAT <= _dmw1_MAT_T_3;
      end
    end
    if (reset) begin
      csrs_28_PLV3 <= 1'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_47) begin
        csrs_28_PLV3 <= rkd[3] & csrMask[3] | csrs_28_PLV3 & ~csrMask[3];
      end
    end
    if (reset) begin
      csrs_28_PLV0 <= 1'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_47) begin
        csrs_28_PLV0 <= _T_1412 | csrs_28_PLV0 & ~csrMask[0];
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_0_E <= _GEN_913;
          end else begin
            tlb_0_E <= _GEN_1939;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_0_VPPN <= _GEN_785;
          end else begin
            tlb_0_VPPN <= _GEN_1811;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_0_PS <= _GEN_817;
          end else begin
            tlb_0_PS <= _GEN_1843;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_0_G <= _GEN_849;
          end else begin
            tlb_0_G <= _GEN_1875;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_0_ASID <= _GEN_881;
          end else begin
            tlb_0_ASID <= _GEN_1907;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_1_E <= _GEN_914;
          end else begin
            tlb_1_E <= _GEN_1940;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_1_VPPN <= _GEN_786;
          end else begin
            tlb_1_VPPN <= _GEN_1812;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_1_PS <= _GEN_818;
          end else begin
            tlb_1_PS <= _GEN_1844;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_1_G <= _GEN_850;
          end else begin
            tlb_1_G <= _GEN_1876;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_1_ASID <= _GEN_882;
          end else begin
            tlb_1_ASID <= _GEN_1908;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_2_E <= _GEN_915;
          end else begin
            tlb_2_E <= _GEN_1941;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_2_VPPN <= _GEN_787;
          end else begin
            tlb_2_VPPN <= _GEN_1813;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_2_PS <= _GEN_819;
          end else begin
            tlb_2_PS <= _GEN_1845;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_2_G <= _GEN_851;
          end else begin
            tlb_2_G <= _GEN_1877;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_2_ASID <= _GEN_883;
          end else begin
            tlb_2_ASID <= _GEN_1909;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_3_E <= _GEN_916;
          end else begin
            tlb_3_E <= _GEN_1942;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_3_VPPN <= _GEN_788;
          end else begin
            tlb_3_VPPN <= _GEN_1814;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_3_PS <= _GEN_820;
          end else begin
            tlb_3_PS <= _GEN_1846;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_3_G <= _GEN_852;
          end else begin
            tlb_3_G <= _GEN_1878;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_3_ASID <= _GEN_884;
          end else begin
            tlb_3_ASID <= _GEN_1910;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_4_E <= _GEN_917;
          end else begin
            tlb_4_E <= _GEN_1943;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_4_VPPN <= _GEN_789;
          end else begin
            tlb_4_VPPN <= _GEN_1815;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_4_PS <= _GEN_821;
          end else begin
            tlb_4_PS <= _GEN_1847;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_4_G <= _GEN_853;
          end else begin
            tlb_4_G <= _GEN_1879;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_4_ASID <= _GEN_885;
          end else begin
            tlb_4_ASID <= _GEN_1911;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_5_E <= _GEN_918;
          end else begin
            tlb_5_E <= _GEN_1944;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_5_VPPN <= _GEN_790;
          end else begin
            tlb_5_VPPN <= _GEN_1816;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_5_PS <= _GEN_822;
          end else begin
            tlb_5_PS <= _GEN_1848;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_5_G <= _GEN_854;
          end else begin
            tlb_5_G <= _GEN_1880;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_5_ASID <= _GEN_886;
          end else begin
            tlb_5_ASID <= _GEN_1912;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_6_E <= _GEN_919;
          end else begin
            tlb_6_E <= _GEN_1945;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_6_VPPN <= _GEN_791;
          end else begin
            tlb_6_VPPN <= _GEN_1817;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_6_PS <= _GEN_823;
          end else begin
            tlb_6_PS <= _GEN_1849;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_6_G <= _GEN_855;
          end else begin
            tlb_6_G <= _GEN_1881;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_6_ASID <= _GEN_887;
          end else begin
            tlb_6_ASID <= _GEN_1913;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_7_E <= _GEN_920;
          end else begin
            tlb_7_E <= _GEN_1946;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_7_VPPN <= _GEN_792;
          end else begin
            tlb_7_VPPN <= _GEN_1818;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_7_PS <= _GEN_824;
          end else begin
            tlb_7_PS <= _GEN_1850;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_7_G <= _GEN_856;
          end else begin
            tlb_7_G <= _GEN_1882;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_7_ASID <= _GEN_888;
          end else begin
            tlb_7_ASID <= _GEN_1914;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_8_E <= _GEN_921;
          end else begin
            tlb_8_E <= _GEN_1947;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_8_VPPN <= _GEN_793;
          end else begin
            tlb_8_VPPN <= _GEN_1819;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_8_PS <= _GEN_825;
          end else begin
            tlb_8_PS <= _GEN_1851;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_8_G <= _GEN_857;
          end else begin
            tlb_8_G <= _GEN_1883;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_8_ASID <= _GEN_889;
          end else begin
            tlb_8_ASID <= _GEN_1915;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_9_E <= _GEN_922;
          end else begin
            tlb_9_E <= _GEN_1948;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_9_VPPN <= _GEN_794;
          end else begin
            tlb_9_VPPN <= _GEN_1820;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_9_PS <= _GEN_826;
          end else begin
            tlb_9_PS <= _GEN_1852;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_9_G <= _GEN_858;
          end else begin
            tlb_9_G <= _GEN_1884;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_9_ASID <= _GEN_890;
          end else begin
            tlb_9_ASID <= _GEN_1916;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_10_E <= _GEN_923;
          end else begin
            tlb_10_E <= _GEN_1949;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_10_VPPN <= _GEN_795;
          end else begin
            tlb_10_VPPN <= _GEN_1821;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_10_PS <= _GEN_827;
          end else begin
            tlb_10_PS <= _GEN_1853;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_10_G <= _GEN_859;
          end else begin
            tlb_10_G <= _GEN_1885;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_10_ASID <= _GEN_891;
          end else begin
            tlb_10_ASID <= _GEN_1917;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_11_E <= _GEN_924;
          end else begin
            tlb_11_E <= _GEN_1950;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_11_VPPN <= _GEN_796;
          end else begin
            tlb_11_VPPN <= _GEN_1822;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_11_PS <= _GEN_828;
          end else begin
            tlb_11_PS <= _GEN_1854;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_11_G <= _GEN_860;
          end else begin
            tlb_11_G <= _GEN_1886;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_11_ASID <= _GEN_892;
          end else begin
            tlb_11_ASID <= _GEN_1918;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_12_E <= _GEN_925;
          end else begin
            tlb_12_E <= _GEN_1951;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_12_VPPN <= _GEN_797;
          end else begin
            tlb_12_VPPN <= _GEN_1823;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_12_PS <= _GEN_829;
          end else begin
            tlb_12_PS <= _GEN_1855;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_12_G <= _GEN_861;
          end else begin
            tlb_12_G <= _GEN_1887;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_12_ASID <= _GEN_893;
          end else begin
            tlb_12_ASID <= _GEN_1919;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_13_E <= _GEN_926;
          end else begin
            tlb_13_E <= _GEN_1952;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_13_VPPN <= _GEN_798;
          end else begin
            tlb_13_VPPN <= _GEN_1824;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_13_PS <= _GEN_830;
          end else begin
            tlb_13_PS <= _GEN_1856;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_13_G <= _GEN_862;
          end else begin
            tlb_13_G <= _GEN_1888;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_13_ASID <= _GEN_894;
          end else begin
            tlb_13_ASID <= _GEN_1920;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_14_E <= _GEN_927;
          end else begin
            tlb_14_E <= _GEN_1953;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_14_VPPN <= _GEN_799;
          end else begin
            tlb_14_VPPN <= _GEN_1825;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_14_PS <= _GEN_831;
          end else begin
            tlb_14_PS <= _GEN_1857;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_14_G <= _GEN_863;
          end else begin
            tlb_14_G <= _GEN_1889;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_14_ASID <= _GEN_895;
          end else begin
            tlb_14_ASID <= _GEN_1921;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_15_E <= _GEN_928;
          end else begin
            tlb_15_E <= _GEN_1954;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_15_VPPN <= _GEN_800;
          end else begin
            tlb_15_VPPN <= _GEN_1826;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_15_PS <= _GEN_832;
          end else begin
            tlb_15_PS <= _GEN_1858;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_15_G <= _GEN_864;
          end else begin
            tlb_15_G <= _GEN_1890;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_15_ASID <= _GEN_896;
          end else begin
            tlb_15_ASID <= _GEN_1922;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_16_E <= _GEN_929;
          end else begin
            tlb_16_E <= _GEN_1955;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_16_VPPN <= _GEN_801;
          end else begin
            tlb_16_VPPN <= _GEN_1827;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_16_PS <= _GEN_833;
          end else begin
            tlb_16_PS <= _GEN_1859;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_16_G <= _GEN_865;
          end else begin
            tlb_16_G <= _GEN_1891;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_16_ASID <= _GEN_897;
          end else begin
            tlb_16_ASID <= _GEN_1923;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_17_E <= _GEN_930;
          end else begin
            tlb_17_E <= _GEN_1956;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_17_VPPN <= _GEN_802;
          end else begin
            tlb_17_VPPN <= _GEN_1828;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_17_PS <= _GEN_834;
          end else begin
            tlb_17_PS <= _GEN_1860;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_17_G <= _GEN_866;
          end else begin
            tlb_17_G <= _GEN_1892;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_17_ASID <= _GEN_898;
          end else begin
            tlb_17_ASID <= _GEN_1924;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_18_E <= _GEN_931;
          end else begin
            tlb_18_E <= _GEN_1957;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_18_VPPN <= _GEN_803;
          end else begin
            tlb_18_VPPN <= _GEN_1829;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_18_PS <= _GEN_835;
          end else begin
            tlb_18_PS <= _GEN_1861;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_18_G <= _GEN_867;
          end else begin
            tlb_18_G <= _GEN_1893;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_18_ASID <= _GEN_899;
          end else begin
            tlb_18_ASID <= _GEN_1925;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_19_E <= _GEN_932;
          end else begin
            tlb_19_E <= _GEN_1958;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_19_VPPN <= _GEN_804;
          end else begin
            tlb_19_VPPN <= _GEN_1830;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_19_PS <= _GEN_836;
          end else begin
            tlb_19_PS <= _GEN_1862;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_19_G <= _GEN_868;
          end else begin
            tlb_19_G <= _GEN_1894;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_19_ASID <= _GEN_900;
          end else begin
            tlb_19_ASID <= _GEN_1926;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_20_E <= _GEN_933;
          end else begin
            tlb_20_E <= _GEN_1959;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_20_VPPN <= _GEN_805;
          end else begin
            tlb_20_VPPN <= _GEN_1831;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_20_PS <= _GEN_837;
          end else begin
            tlb_20_PS <= _GEN_1863;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_20_G <= _GEN_869;
          end else begin
            tlb_20_G <= _GEN_1895;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_20_ASID <= _GEN_901;
          end else begin
            tlb_20_ASID <= _GEN_1927;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_21_E <= _GEN_934;
          end else begin
            tlb_21_E <= _GEN_1960;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_21_VPPN <= _GEN_806;
          end else begin
            tlb_21_VPPN <= _GEN_1832;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_21_PS <= _GEN_838;
          end else begin
            tlb_21_PS <= _GEN_1864;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_21_G <= _GEN_870;
          end else begin
            tlb_21_G <= _GEN_1896;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_21_ASID <= _GEN_902;
          end else begin
            tlb_21_ASID <= _GEN_1928;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_22_E <= _GEN_935;
          end else begin
            tlb_22_E <= _GEN_1961;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_22_VPPN <= _GEN_807;
          end else begin
            tlb_22_VPPN <= _GEN_1833;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_22_PS <= _GEN_839;
          end else begin
            tlb_22_PS <= _GEN_1865;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_22_G <= _GEN_871;
          end else begin
            tlb_22_G <= _GEN_1897;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_22_ASID <= _GEN_903;
          end else begin
            tlb_22_ASID <= _GEN_1929;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_23_E <= _GEN_936;
          end else begin
            tlb_23_E <= _GEN_1962;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_23_VPPN <= _GEN_808;
          end else begin
            tlb_23_VPPN <= _GEN_1834;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_23_PS <= _GEN_840;
          end else begin
            tlb_23_PS <= _GEN_1866;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_23_G <= _GEN_872;
          end else begin
            tlb_23_G <= _GEN_1898;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_23_ASID <= _GEN_904;
          end else begin
            tlb_23_ASID <= _GEN_1930;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_24_E <= _GEN_937;
          end else begin
            tlb_24_E <= _GEN_1963;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_24_VPPN <= _GEN_809;
          end else begin
            tlb_24_VPPN <= _GEN_1835;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_24_PS <= _GEN_841;
          end else begin
            tlb_24_PS <= _GEN_1867;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_24_G <= _GEN_873;
          end else begin
            tlb_24_G <= _GEN_1899;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_24_ASID <= _GEN_905;
          end else begin
            tlb_24_ASID <= _GEN_1931;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_25_E <= _GEN_938;
          end else begin
            tlb_25_E <= _GEN_1964;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_25_VPPN <= _GEN_810;
          end else begin
            tlb_25_VPPN <= _GEN_1836;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_25_PS <= _GEN_842;
          end else begin
            tlb_25_PS <= _GEN_1868;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_25_G <= _GEN_874;
          end else begin
            tlb_25_G <= _GEN_1900;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_25_ASID <= _GEN_906;
          end else begin
            tlb_25_ASID <= _GEN_1932;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_26_E <= _GEN_939;
          end else begin
            tlb_26_E <= _GEN_1965;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_26_VPPN <= _GEN_811;
          end else begin
            tlb_26_VPPN <= _GEN_1837;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_26_PS <= _GEN_843;
          end else begin
            tlb_26_PS <= _GEN_1869;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_26_G <= _GEN_875;
          end else begin
            tlb_26_G <= _GEN_1901;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_26_ASID <= _GEN_907;
          end else begin
            tlb_26_ASID <= _GEN_1933;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_27_E <= _GEN_940;
          end else begin
            tlb_27_E <= _GEN_1966;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_27_VPPN <= _GEN_812;
          end else begin
            tlb_27_VPPN <= _GEN_1838;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_27_PS <= _GEN_844;
          end else begin
            tlb_27_PS <= _GEN_1870;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_27_G <= _GEN_876;
          end else begin
            tlb_27_G <= _GEN_1902;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_27_ASID <= _GEN_908;
          end else begin
            tlb_27_ASID <= _GEN_1934;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_28_E <= _GEN_941;
          end else begin
            tlb_28_E <= _GEN_1967;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_28_VPPN <= _GEN_813;
          end else begin
            tlb_28_VPPN <= _GEN_1839;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_28_PS <= _GEN_845;
          end else begin
            tlb_28_PS <= _GEN_1871;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_28_G <= _GEN_877;
          end else begin
            tlb_28_G <= _GEN_1903;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_28_ASID <= _GEN_909;
          end else begin
            tlb_28_ASID <= _GEN_1935;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_29_E <= _GEN_942;
          end else begin
            tlb_29_E <= _GEN_1968;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_29_VPPN <= _GEN_814;
          end else begin
            tlb_29_VPPN <= _GEN_1840;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_29_PS <= _GEN_846;
          end else begin
            tlb_29_PS <= _GEN_1872;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_29_G <= _GEN_878;
          end else begin
            tlb_29_G <= _GEN_1904;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_29_ASID <= _GEN_910;
          end else begin
            tlb_29_ASID <= _GEN_1936;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_30_E <= _GEN_943;
          end else begin
            tlb_30_E <= _GEN_1969;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_30_VPPN <= _GEN_815;
          end else begin
            tlb_30_VPPN <= _GEN_1841;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_30_PS <= _GEN_847;
          end else begin
            tlb_30_PS <= _GEN_1873;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_30_G <= _GEN_879;
          end else begin
            tlb_30_G <= _GEN_1905;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_30_ASID <= _GEN_911;
          end else begin
            tlb_30_ASID <= _GEN_1937;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_31_E <= _GEN_944;
          end else begin
            tlb_31_E <= _GEN_1970;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_31_VPPN <= _GEN_816;
          end else begin
            tlb_31_VPPN <= _GEN_1842;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_31_PS <= _GEN_848;
          end else begin
            tlb_31_PS <= _GEN_1874;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_31_G <= _GEN_880;
          end else begin
            tlb_31_G <= _GEN_1906;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_31_ASID <= _GEN_912;
          end else begin
            tlb_31_ASID <= _GEN_1938;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_0_P1_V <= _GEN_1233;
          end else begin
            tlb_0_P1_V <= _GEN_2259;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_1_P1_V <= _GEN_1234;
          end else begin
            tlb_1_P1_V <= _GEN_2260;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_2_P1_V <= _GEN_1235;
          end else begin
            tlb_2_P1_V <= _GEN_2261;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_3_P1_V <= _GEN_1236;
          end else begin
            tlb_3_P1_V <= _GEN_2262;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_4_P1_V <= _GEN_1237;
          end else begin
            tlb_4_P1_V <= _GEN_2263;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_5_P1_V <= _GEN_1238;
          end else begin
            tlb_5_P1_V <= _GEN_2264;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_6_P1_V <= _GEN_1239;
          end else begin
            tlb_6_P1_V <= _GEN_2265;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_7_P1_V <= _GEN_1240;
          end else begin
            tlb_7_P1_V <= _GEN_2266;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_8_P1_V <= _GEN_1241;
          end else begin
            tlb_8_P1_V <= _GEN_2267;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_9_P1_V <= _GEN_1242;
          end else begin
            tlb_9_P1_V <= _GEN_2268;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_10_P1_V <= _GEN_1243;
          end else begin
            tlb_10_P1_V <= _GEN_2269;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_11_P1_V <= _GEN_1244;
          end else begin
            tlb_11_P1_V <= _GEN_2270;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_12_P1_V <= _GEN_1245;
          end else begin
            tlb_12_P1_V <= _GEN_2271;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_13_P1_V <= _GEN_1246;
          end else begin
            tlb_13_P1_V <= _GEN_2272;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_14_P1_V <= _GEN_1247;
          end else begin
            tlb_14_P1_V <= _GEN_2273;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_15_P1_V <= _GEN_1248;
          end else begin
            tlb_15_P1_V <= _GEN_2274;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_16_P1_V <= _GEN_1249;
          end else begin
            tlb_16_P1_V <= _GEN_2275;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_17_P1_V <= _GEN_1250;
          end else begin
            tlb_17_P1_V <= _GEN_2276;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_18_P1_V <= _GEN_1251;
          end else begin
            tlb_18_P1_V <= _GEN_2277;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_19_P1_V <= _GEN_1252;
          end else begin
            tlb_19_P1_V <= _GEN_2278;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_20_P1_V <= _GEN_1253;
          end else begin
            tlb_20_P1_V <= _GEN_2279;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_21_P1_V <= _GEN_1254;
          end else begin
            tlb_21_P1_V <= _GEN_2280;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_22_P1_V <= _GEN_1255;
          end else begin
            tlb_22_P1_V <= _GEN_2281;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_23_P1_V <= _GEN_1256;
          end else begin
            tlb_23_P1_V <= _GEN_2282;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_24_P1_V <= _GEN_1257;
          end else begin
            tlb_24_P1_V <= _GEN_2283;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_25_P1_V <= _GEN_1258;
          end else begin
            tlb_25_P1_V <= _GEN_2284;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_26_P1_V <= _GEN_1259;
          end else begin
            tlb_26_P1_V <= _GEN_2285;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_27_P1_V <= _GEN_1260;
          end else begin
            tlb_27_P1_V <= _GEN_2286;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_28_P1_V <= _GEN_1261;
          end else begin
            tlb_28_P1_V <= _GEN_2287;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_29_P1_V <= _GEN_1262;
          end else begin
            tlb_29_P1_V <= _GEN_2288;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_30_P1_V <= _GEN_1263;
          end else begin
            tlb_30_P1_V <= _GEN_2289;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_31_P1_V <= _GEN_1264;
          end else begin
            tlb_31_P1_V <= _GEN_2290;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_0_P0_V <= _GEN_1073;
          end else begin
            tlb_0_P0_V <= _GEN_2099;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_1_P0_V <= _GEN_1074;
          end else begin
            tlb_1_P0_V <= _GEN_2100;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_2_P0_V <= _GEN_1075;
          end else begin
            tlb_2_P0_V <= _GEN_2101;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_3_P0_V <= _GEN_1076;
          end else begin
            tlb_3_P0_V <= _GEN_2102;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_4_P0_V <= _GEN_1077;
          end else begin
            tlb_4_P0_V <= _GEN_2103;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_5_P0_V <= _GEN_1078;
          end else begin
            tlb_5_P0_V <= _GEN_2104;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_6_P0_V <= _GEN_1079;
          end else begin
            tlb_6_P0_V <= _GEN_2105;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_7_P0_V <= _GEN_1080;
          end else begin
            tlb_7_P0_V <= _GEN_2106;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_8_P0_V <= _GEN_1081;
          end else begin
            tlb_8_P0_V <= _GEN_2107;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_9_P0_V <= _GEN_1082;
          end else begin
            tlb_9_P0_V <= _GEN_2108;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_10_P0_V <= _GEN_1083;
          end else begin
            tlb_10_P0_V <= _GEN_2109;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_11_P0_V <= _GEN_1084;
          end else begin
            tlb_11_P0_V <= _GEN_2110;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_12_P0_V <= _GEN_1085;
          end else begin
            tlb_12_P0_V <= _GEN_2111;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_13_P0_V <= _GEN_1086;
          end else begin
            tlb_13_P0_V <= _GEN_2112;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_14_P0_V <= _GEN_1087;
          end else begin
            tlb_14_P0_V <= _GEN_2113;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_15_P0_V <= _GEN_1088;
          end else begin
            tlb_15_P0_V <= _GEN_2114;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_16_P0_V <= _GEN_1089;
          end else begin
            tlb_16_P0_V <= _GEN_2115;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_17_P0_V <= _GEN_1090;
          end else begin
            tlb_17_P0_V <= _GEN_2116;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_18_P0_V <= _GEN_1091;
          end else begin
            tlb_18_P0_V <= _GEN_2117;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_19_P0_V <= _GEN_1092;
          end else begin
            tlb_19_P0_V <= _GEN_2118;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_20_P0_V <= _GEN_1093;
          end else begin
            tlb_20_P0_V <= _GEN_2119;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_21_P0_V <= _GEN_1094;
          end else begin
            tlb_21_P0_V <= _GEN_2120;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_22_P0_V <= _GEN_1095;
          end else begin
            tlb_22_P0_V <= _GEN_2121;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_23_P0_V <= _GEN_1096;
          end else begin
            tlb_23_P0_V <= _GEN_2122;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_24_P0_V <= _GEN_1097;
          end else begin
            tlb_24_P0_V <= _GEN_2123;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_25_P0_V <= _GEN_1098;
          end else begin
            tlb_25_P0_V <= _GEN_2124;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_26_P0_V <= _GEN_1099;
          end else begin
            tlb_26_P0_V <= _GEN_2125;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_27_P0_V <= _GEN_1100;
          end else begin
            tlb_27_P0_V <= _GEN_2126;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_28_P0_V <= _GEN_1101;
          end else begin
            tlb_28_P0_V <= _GEN_2127;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_29_P0_V <= _GEN_1102;
          end else begin
            tlb_29_P0_V <= _GEN_2128;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_30_P0_V <= _GEN_1103;
          end else begin
            tlb_30_P0_V <= _GEN_2129;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_31_P0_V <= _GEN_1104;
          end else begin
            tlb_31_P0_V <= _GEN_2130;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_0_P1_PLV <= _GEN_1137;
          end else begin
            tlb_0_P1_PLV <= _GEN_2163;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_1_P1_PLV <= _GEN_1138;
          end else begin
            tlb_1_P1_PLV <= _GEN_2164;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_2_P1_PLV <= _GEN_1139;
          end else begin
            tlb_2_P1_PLV <= _GEN_2165;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_3_P1_PLV <= _GEN_1140;
          end else begin
            tlb_3_P1_PLV <= _GEN_2166;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_4_P1_PLV <= _GEN_1141;
          end else begin
            tlb_4_P1_PLV <= _GEN_2167;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_5_P1_PLV <= _GEN_1142;
          end else begin
            tlb_5_P1_PLV <= _GEN_2168;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_6_P1_PLV <= _GEN_1143;
          end else begin
            tlb_6_P1_PLV <= _GEN_2169;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_7_P1_PLV <= _GEN_1144;
          end else begin
            tlb_7_P1_PLV <= _GEN_2170;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_8_P1_PLV <= _GEN_1145;
          end else begin
            tlb_8_P1_PLV <= _GEN_2171;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_9_P1_PLV <= _GEN_1146;
          end else begin
            tlb_9_P1_PLV <= _GEN_2172;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_10_P1_PLV <= _GEN_1147;
          end else begin
            tlb_10_P1_PLV <= _GEN_2173;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_11_P1_PLV <= _GEN_1148;
          end else begin
            tlb_11_P1_PLV <= _GEN_2174;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_12_P1_PLV <= _GEN_1149;
          end else begin
            tlb_12_P1_PLV <= _GEN_2175;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_13_P1_PLV <= _GEN_1150;
          end else begin
            tlb_13_P1_PLV <= _GEN_2176;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_14_P1_PLV <= _GEN_1151;
          end else begin
            tlb_14_P1_PLV <= _GEN_2177;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_15_P1_PLV <= _GEN_1152;
          end else begin
            tlb_15_P1_PLV <= _GEN_2178;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_16_P1_PLV <= _GEN_1153;
          end else begin
            tlb_16_P1_PLV <= _GEN_2179;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_17_P1_PLV <= _GEN_1154;
          end else begin
            tlb_17_P1_PLV <= _GEN_2180;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_18_P1_PLV <= _GEN_1155;
          end else begin
            tlb_18_P1_PLV <= _GEN_2181;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_19_P1_PLV <= _GEN_1156;
          end else begin
            tlb_19_P1_PLV <= _GEN_2182;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_20_P1_PLV <= _GEN_1157;
          end else begin
            tlb_20_P1_PLV <= _GEN_2183;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_21_P1_PLV <= _GEN_1158;
          end else begin
            tlb_21_P1_PLV <= _GEN_2184;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_22_P1_PLV <= _GEN_1159;
          end else begin
            tlb_22_P1_PLV <= _GEN_2185;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_23_P1_PLV <= _GEN_1160;
          end else begin
            tlb_23_P1_PLV <= _GEN_2186;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_24_P1_PLV <= _GEN_1161;
          end else begin
            tlb_24_P1_PLV <= _GEN_2187;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_25_P1_PLV <= _GEN_1162;
          end else begin
            tlb_25_P1_PLV <= _GEN_2188;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_26_P1_PLV <= _GEN_1163;
          end else begin
            tlb_26_P1_PLV <= _GEN_2189;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_27_P1_PLV <= _GEN_1164;
          end else begin
            tlb_27_P1_PLV <= _GEN_2190;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_28_P1_PLV <= _GEN_1165;
          end else begin
            tlb_28_P1_PLV <= _GEN_2191;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_29_P1_PLV <= _GEN_1166;
          end else begin
            tlb_29_P1_PLV <= _GEN_2192;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_30_P1_PLV <= _GEN_1167;
          end else begin
            tlb_30_P1_PLV <= _GEN_2193;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_31_P1_PLV <= _GEN_1168;
          end else begin
            tlb_31_P1_PLV <= _GEN_2194;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_0_P0_PLV <= _GEN_977;
          end else begin
            tlb_0_P0_PLV <= _GEN_2003;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_1_P0_PLV <= _GEN_978;
          end else begin
            tlb_1_P0_PLV <= _GEN_2004;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_2_P0_PLV <= _GEN_979;
          end else begin
            tlb_2_P0_PLV <= _GEN_2005;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_3_P0_PLV <= _GEN_980;
          end else begin
            tlb_3_P0_PLV <= _GEN_2006;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_4_P0_PLV <= _GEN_981;
          end else begin
            tlb_4_P0_PLV <= _GEN_2007;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_5_P0_PLV <= _GEN_982;
          end else begin
            tlb_5_P0_PLV <= _GEN_2008;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_6_P0_PLV <= _GEN_983;
          end else begin
            tlb_6_P0_PLV <= _GEN_2009;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_7_P0_PLV <= _GEN_984;
          end else begin
            tlb_7_P0_PLV <= _GEN_2010;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_8_P0_PLV <= _GEN_985;
          end else begin
            tlb_8_P0_PLV <= _GEN_2011;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_9_P0_PLV <= _GEN_986;
          end else begin
            tlb_9_P0_PLV <= _GEN_2012;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_10_P0_PLV <= _GEN_987;
          end else begin
            tlb_10_P0_PLV <= _GEN_2013;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_11_P0_PLV <= _GEN_988;
          end else begin
            tlb_11_P0_PLV <= _GEN_2014;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_12_P0_PLV <= _GEN_989;
          end else begin
            tlb_12_P0_PLV <= _GEN_2015;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_13_P0_PLV <= _GEN_990;
          end else begin
            tlb_13_P0_PLV <= _GEN_2016;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_14_P0_PLV <= _GEN_991;
          end else begin
            tlb_14_P0_PLV <= _GEN_2017;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_15_P0_PLV <= _GEN_992;
          end else begin
            tlb_15_P0_PLV <= _GEN_2018;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_16_P0_PLV <= _GEN_993;
          end else begin
            tlb_16_P0_PLV <= _GEN_2019;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_17_P0_PLV <= _GEN_994;
          end else begin
            tlb_17_P0_PLV <= _GEN_2020;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_18_P0_PLV <= _GEN_995;
          end else begin
            tlb_18_P0_PLV <= _GEN_2021;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_19_P0_PLV <= _GEN_996;
          end else begin
            tlb_19_P0_PLV <= _GEN_2022;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_20_P0_PLV <= _GEN_997;
          end else begin
            tlb_20_P0_PLV <= _GEN_2023;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_21_P0_PLV <= _GEN_998;
          end else begin
            tlb_21_P0_PLV <= _GEN_2024;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_22_P0_PLV <= _GEN_999;
          end else begin
            tlb_22_P0_PLV <= _GEN_2025;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_23_P0_PLV <= _GEN_1000;
          end else begin
            tlb_23_P0_PLV <= _GEN_2026;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_24_P0_PLV <= _GEN_1001;
          end else begin
            tlb_24_P0_PLV <= _GEN_2027;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_25_P0_PLV <= _GEN_1002;
          end else begin
            tlb_25_P0_PLV <= _GEN_2028;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_26_P0_PLV <= _GEN_1003;
          end else begin
            tlb_26_P0_PLV <= _GEN_2029;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_27_P0_PLV <= _GEN_1004;
          end else begin
            tlb_27_P0_PLV <= _GEN_2030;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_28_P0_PLV <= _GEN_1005;
          end else begin
            tlb_28_P0_PLV <= _GEN_2031;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_29_P0_PLV <= _GEN_1006;
          end else begin
            tlb_29_P0_PLV <= _GEN_2032;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_30_P0_PLV <= _GEN_1007;
          end else begin
            tlb_30_P0_PLV <= _GEN_2033;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_31_P0_PLV <= _GEN_1008;
          end else begin
            tlb_31_P0_PLV <= _GEN_2034;
          end
        end
      end
    end
    if (!(dStallReg)) begin
      inst_reg <= io_inst_resp_bits;
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_0_P1_D <= _GEN_1201;
          end else begin
            tlb_0_P1_D <= _GEN_2227;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_1_P1_D <= _GEN_1202;
          end else begin
            tlb_1_P1_D <= _GEN_2228;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_2_P1_D <= _GEN_1203;
          end else begin
            tlb_2_P1_D <= _GEN_2229;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_3_P1_D <= _GEN_1204;
          end else begin
            tlb_3_P1_D <= _GEN_2230;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_4_P1_D <= _GEN_1205;
          end else begin
            tlb_4_P1_D <= _GEN_2231;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_5_P1_D <= _GEN_1206;
          end else begin
            tlb_5_P1_D <= _GEN_2232;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_6_P1_D <= _GEN_1207;
          end else begin
            tlb_6_P1_D <= _GEN_2233;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_7_P1_D <= _GEN_1208;
          end else begin
            tlb_7_P1_D <= _GEN_2234;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_8_P1_D <= _GEN_1209;
          end else begin
            tlb_8_P1_D <= _GEN_2235;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_9_P1_D <= _GEN_1210;
          end else begin
            tlb_9_P1_D <= _GEN_2236;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_10_P1_D <= _GEN_1211;
          end else begin
            tlb_10_P1_D <= _GEN_2237;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_11_P1_D <= _GEN_1212;
          end else begin
            tlb_11_P1_D <= _GEN_2238;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_12_P1_D <= _GEN_1213;
          end else begin
            tlb_12_P1_D <= _GEN_2239;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_13_P1_D <= _GEN_1214;
          end else begin
            tlb_13_P1_D <= _GEN_2240;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_14_P1_D <= _GEN_1215;
          end else begin
            tlb_14_P1_D <= _GEN_2241;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_15_P1_D <= _GEN_1216;
          end else begin
            tlb_15_P1_D <= _GEN_2242;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_16_P1_D <= _GEN_1217;
          end else begin
            tlb_16_P1_D <= _GEN_2243;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_17_P1_D <= _GEN_1218;
          end else begin
            tlb_17_P1_D <= _GEN_2244;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_18_P1_D <= _GEN_1219;
          end else begin
            tlb_18_P1_D <= _GEN_2245;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_19_P1_D <= _GEN_1220;
          end else begin
            tlb_19_P1_D <= _GEN_2246;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_20_P1_D <= _GEN_1221;
          end else begin
            tlb_20_P1_D <= _GEN_2247;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_21_P1_D <= _GEN_1222;
          end else begin
            tlb_21_P1_D <= _GEN_2248;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_22_P1_D <= _GEN_1223;
          end else begin
            tlb_22_P1_D <= _GEN_2249;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_23_P1_D <= _GEN_1224;
          end else begin
            tlb_23_P1_D <= _GEN_2250;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_24_P1_D <= _GEN_1225;
          end else begin
            tlb_24_P1_D <= _GEN_2251;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_25_P1_D <= _GEN_1226;
          end else begin
            tlb_25_P1_D <= _GEN_2252;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_26_P1_D <= _GEN_1227;
          end else begin
            tlb_26_P1_D <= _GEN_2253;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_27_P1_D <= _GEN_1228;
          end else begin
            tlb_27_P1_D <= _GEN_2254;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_28_P1_D <= _GEN_1229;
          end else begin
            tlb_28_P1_D <= _GEN_2255;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_29_P1_D <= _GEN_1230;
          end else begin
            tlb_29_P1_D <= _GEN_2256;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_30_P1_D <= _GEN_1231;
          end else begin
            tlb_30_P1_D <= _GEN_2257;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_31_P1_D <= _GEN_1232;
          end else begin
            tlb_31_P1_D <= _GEN_2258;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_0_P0_D <= _GEN_1041;
          end else begin
            tlb_0_P0_D <= _GEN_2067;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_1_P0_D <= _GEN_1042;
          end else begin
            tlb_1_P0_D <= _GEN_2068;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_2_P0_D <= _GEN_1043;
          end else begin
            tlb_2_P0_D <= _GEN_2069;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_3_P0_D <= _GEN_1044;
          end else begin
            tlb_3_P0_D <= _GEN_2070;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_4_P0_D <= _GEN_1045;
          end else begin
            tlb_4_P0_D <= _GEN_2071;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_5_P0_D <= _GEN_1046;
          end else begin
            tlb_5_P0_D <= _GEN_2072;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_6_P0_D <= _GEN_1047;
          end else begin
            tlb_6_P0_D <= _GEN_2073;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_7_P0_D <= _GEN_1048;
          end else begin
            tlb_7_P0_D <= _GEN_2074;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_8_P0_D <= _GEN_1049;
          end else begin
            tlb_8_P0_D <= _GEN_2075;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_9_P0_D <= _GEN_1050;
          end else begin
            tlb_9_P0_D <= _GEN_2076;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_10_P0_D <= _GEN_1051;
          end else begin
            tlb_10_P0_D <= _GEN_2077;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_11_P0_D <= _GEN_1052;
          end else begin
            tlb_11_P0_D <= _GEN_2078;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_12_P0_D <= _GEN_1053;
          end else begin
            tlb_12_P0_D <= _GEN_2079;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_13_P0_D <= _GEN_1054;
          end else begin
            tlb_13_P0_D <= _GEN_2080;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_14_P0_D <= _GEN_1055;
          end else begin
            tlb_14_P0_D <= _GEN_2081;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_15_P0_D <= _GEN_1056;
          end else begin
            tlb_15_P0_D <= _GEN_2082;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_16_P0_D <= _GEN_1057;
          end else begin
            tlb_16_P0_D <= _GEN_2083;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_17_P0_D <= _GEN_1058;
          end else begin
            tlb_17_P0_D <= _GEN_2084;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_18_P0_D <= _GEN_1059;
          end else begin
            tlb_18_P0_D <= _GEN_2085;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_19_P0_D <= _GEN_1060;
          end else begin
            tlb_19_P0_D <= _GEN_2086;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_20_P0_D <= _GEN_1061;
          end else begin
            tlb_20_P0_D <= _GEN_2087;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_21_P0_D <= _GEN_1062;
          end else begin
            tlb_21_P0_D <= _GEN_2088;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_22_P0_D <= _GEN_1063;
          end else begin
            tlb_22_P0_D <= _GEN_2089;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_23_P0_D <= _GEN_1064;
          end else begin
            tlb_23_P0_D <= _GEN_2090;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_24_P0_D <= _GEN_1065;
          end else begin
            tlb_24_P0_D <= _GEN_2091;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_25_P0_D <= _GEN_1066;
          end else begin
            tlb_25_P0_D <= _GEN_2092;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_26_P0_D <= _GEN_1067;
          end else begin
            tlb_26_P0_D <= _GEN_2093;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_27_P0_D <= _GEN_1068;
          end else begin
            tlb_27_P0_D <= _GEN_2094;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_28_P0_D <= _GEN_1069;
          end else begin
            tlb_28_P0_D <= _GEN_2095;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_29_P0_D <= _GEN_1070;
          end else begin
            tlb_29_P0_D <= _GEN_2096;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_30_P0_D <= _GEN_1071;
          end else begin
            tlb_30_P0_D <= _GEN_2097;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_31_P0_D <= _GEN_1072;
          end else begin
            tlb_31_P0_D <= _GEN_2098;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_0_P0_PPN <= _GEN_945;
          end else begin
            tlb_0_P0_PPN <= _GEN_1971;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_0_P0_MAT <= _GEN_1009;
          end else begin
            tlb_0_P0_MAT <= _GEN_2035;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_0_P1_PPN <= _GEN_1105;
          end else begin
            tlb_0_P1_PPN <= _GEN_2131;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_0_P1_MAT <= _GEN_1169;
          end else begin
            tlb_0_P1_MAT <= _GEN_2195;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_1_P0_PPN <= _GEN_946;
          end else begin
            tlb_1_P0_PPN <= _GEN_1972;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_1_P0_MAT <= _GEN_1010;
          end else begin
            tlb_1_P0_MAT <= _GEN_2036;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_1_P1_PPN <= _GEN_1106;
          end else begin
            tlb_1_P1_PPN <= _GEN_2132;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_1_P1_MAT <= _GEN_1170;
          end else begin
            tlb_1_P1_MAT <= _GEN_2196;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_2_P0_PPN <= _GEN_947;
          end else begin
            tlb_2_P0_PPN <= _GEN_1973;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_2_P0_MAT <= _GEN_1011;
          end else begin
            tlb_2_P0_MAT <= _GEN_2037;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_2_P1_PPN <= _GEN_1107;
          end else begin
            tlb_2_P1_PPN <= _GEN_2133;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_2_P1_MAT <= _GEN_1171;
          end else begin
            tlb_2_P1_MAT <= _GEN_2197;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_3_P0_PPN <= _GEN_948;
          end else begin
            tlb_3_P0_PPN <= _GEN_1974;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_3_P0_MAT <= _GEN_1012;
          end else begin
            tlb_3_P0_MAT <= _GEN_2038;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_3_P1_PPN <= _GEN_1108;
          end else begin
            tlb_3_P1_PPN <= _GEN_2134;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_3_P1_MAT <= _GEN_1172;
          end else begin
            tlb_3_P1_MAT <= _GEN_2198;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_4_P0_PPN <= _GEN_949;
          end else begin
            tlb_4_P0_PPN <= _GEN_1975;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_4_P0_MAT <= _GEN_1013;
          end else begin
            tlb_4_P0_MAT <= _GEN_2039;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_4_P1_PPN <= _GEN_1109;
          end else begin
            tlb_4_P1_PPN <= _GEN_2135;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_4_P1_MAT <= _GEN_1173;
          end else begin
            tlb_4_P1_MAT <= _GEN_2199;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_5_P0_PPN <= _GEN_950;
          end else begin
            tlb_5_P0_PPN <= _GEN_1976;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_5_P0_MAT <= _GEN_1014;
          end else begin
            tlb_5_P0_MAT <= _GEN_2040;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_5_P1_PPN <= _GEN_1110;
          end else begin
            tlb_5_P1_PPN <= _GEN_2136;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_5_P1_MAT <= _GEN_1174;
          end else begin
            tlb_5_P1_MAT <= _GEN_2200;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_6_P0_PPN <= _GEN_951;
          end else begin
            tlb_6_P0_PPN <= _GEN_1977;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_6_P0_MAT <= _GEN_1015;
          end else begin
            tlb_6_P0_MAT <= _GEN_2041;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_6_P1_PPN <= _GEN_1111;
          end else begin
            tlb_6_P1_PPN <= _GEN_2137;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_6_P1_MAT <= _GEN_1175;
          end else begin
            tlb_6_P1_MAT <= _GEN_2201;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_7_P0_PPN <= _GEN_952;
          end else begin
            tlb_7_P0_PPN <= _GEN_1978;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_7_P0_MAT <= _GEN_1016;
          end else begin
            tlb_7_P0_MAT <= _GEN_2042;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_7_P1_PPN <= _GEN_1112;
          end else begin
            tlb_7_P1_PPN <= _GEN_2138;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_7_P1_MAT <= _GEN_1176;
          end else begin
            tlb_7_P1_MAT <= _GEN_2202;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_8_P0_PPN <= _GEN_953;
          end else begin
            tlb_8_P0_PPN <= _GEN_1979;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_8_P0_MAT <= _GEN_1017;
          end else begin
            tlb_8_P0_MAT <= _GEN_2043;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_8_P1_PPN <= _GEN_1113;
          end else begin
            tlb_8_P1_PPN <= _GEN_2139;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_8_P1_MAT <= _GEN_1177;
          end else begin
            tlb_8_P1_MAT <= _GEN_2203;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_9_P0_PPN <= _GEN_954;
          end else begin
            tlb_9_P0_PPN <= _GEN_1980;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_9_P0_MAT <= _GEN_1018;
          end else begin
            tlb_9_P0_MAT <= _GEN_2044;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_9_P1_PPN <= _GEN_1114;
          end else begin
            tlb_9_P1_PPN <= _GEN_2140;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_9_P1_MAT <= _GEN_1178;
          end else begin
            tlb_9_P1_MAT <= _GEN_2204;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_10_P0_PPN <= _GEN_955;
          end else begin
            tlb_10_P0_PPN <= _GEN_1981;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_10_P0_MAT <= _GEN_1019;
          end else begin
            tlb_10_P0_MAT <= _GEN_2045;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_10_P1_PPN <= _GEN_1115;
          end else begin
            tlb_10_P1_PPN <= _GEN_2141;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_10_P1_MAT <= _GEN_1179;
          end else begin
            tlb_10_P1_MAT <= _GEN_2205;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_11_P0_PPN <= _GEN_956;
          end else begin
            tlb_11_P0_PPN <= _GEN_1982;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_11_P0_MAT <= _GEN_1020;
          end else begin
            tlb_11_P0_MAT <= _GEN_2046;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_11_P1_PPN <= _GEN_1116;
          end else begin
            tlb_11_P1_PPN <= _GEN_2142;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_11_P1_MAT <= _GEN_1180;
          end else begin
            tlb_11_P1_MAT <= _GEN_2206;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_12_P0_PPN <= _GEN_957;
          end else begin
            tlb_12_P0_PPN <= _GEN_1983;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_12_P0_MAT <= _GEN_1021;
          end else begin
            tlb_12_P0_MAT <= _GEN_2047;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_12_P1_PPN <= _GEN_1117;
          end else begin
            tlb_12_P1_PPN <= _GEN_2143;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_12_P1_MAT <= _GEN_1181;
          end else begin
            tlb_12_P1_MAT <= _GEN_2207;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_13_P0_PPN <= _GEN_958;
          end else begin
            tlb_13_P0_PPN <= _GEN_1984;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_13_P0_MAT <= _GEN_1022;
          end else begin
            tlb_13_P0_MAT <= _GEN_2048;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_13_P1_PPN <= _GEN_1118;
          end else begin
            tlb_13_P1_PPN <= _GEN_2144;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_13_P1_MAT <= _GEN_1182;
          end else begin
            tlb_13_P1_MAT <= _GEN_2208;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_14_P0_PPN <= _GEN_959;
          end else begin
            tlb_14_P0_PPN <= _GEN_1985;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_14_P0_MAT <= _GEN_1023;
          end else begin
            tlb_14_P0_MAT <= _GEN_2049;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_14_P1_PPN <= _GEN_1119;
          end else begin
            tlb_14_P1_PPN <= _GEN_2145;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_14_P1_MAT <= _GEN_1183;
          end else begin
            tlb_14_P1_MAT <= _GEN_2209;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_15_P0_PPN <= _GEN_960;
          end else begin
            tlb_15_P0_PPN <= _GEN_1986;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_15_P0_MAT <= _GEN_1024;
          end else begin
            tlb_15_P0_MAT <= _GEN_2050;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_15_P1_PPN <= _GEN_1120;
          end else begin
            tlb_15_P1_PPN <= _GEN_2146;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_15_P1_MAT <= _GEN_1184;
          end else begin
            tlb_15_P1_MAT <= _GEN_2210;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_16_P0_PPN <= _GEN_961;
          end else begin
            tlb_16_P0_PPN <= _GEN_1987;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_16_P0_MAT <= _GEN_1025;
          end else begin
            tlb_16_P0_MAT <= _GEN_2051;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_16_P1_PPN <= _GEN_1121;
          end else begin
            tlb_16_P1_PPN <= _GEN_2147;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_16_P1_MAT <= _GEN_1185;
          end else begin
            tlb_16_P1_MAT <= _GEN_2211;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_17_P0_PPN <= _GEN_962;
          end else begin
            tlb_17_P0_PPN <= _GEN_1988;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_17_P0_MAT <= _GEN_1026;
          end else begin
            tlb_17_P0_MAT <= _GEN_2052;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_17_P1_PPN <= _GEN_1122;
          end else begin
            tlb_17_P1_PPN <= _GEN_2148;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_17_P1_MAT <= _GEN_1186;
          end else begin
            tlb_17_P1_MAT <= _GEN_2212;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_18_P0_PPN <= _GEN_963;
          end else begin
            tlb_18_P0_PPN <= _GEN_1989;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_18_P0_MAT <= _GEN_1027;
          end else begin
            tlb_18_P0_MAT <= _GEN_2053;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_18_P1_PPN <= _GEN_1123;
          end else begin
            tlb_18_P1_PPN <= _GEN_2149;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_18_P1_MAT <= _GEN_1187;
          end else begin
            tlb_18_P1_MAT <= _GEN_2213;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_19_P0_PPN <= _GEN_964;
          end else begin
            tlb_19_P0_PPN <= _GEN_1990;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_19_P0_MAT <= _GEN_1028;
          end else begin
            tlb_19_P0_MAT <= _GEN_2054;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_19_P1_PPN <= _GEN_1124;
          end else begin
            tlb_19_P1_PPN <= _GEN_2150;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_19_P1_MAT <= _GEN_1188;
          end else begin
            tlb_19_P1_MAT <= _GEN_2214;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_20_P0_PPN <= _GEN_965;
          end else begin
            tlb_20_P0_PPN <= _GEN_1991;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_20_P0_MAT <= _GEN_1029;
          end else begin
            tlb_20_P0_MAT <= _GEN_2055;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_20_P1_PPN <= _GEN_1125;
          end else begin
            tlb_20_P1_PPN <= _GEN_2151;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_20_P1_MAT <= _GEN_1189;
          end else begin
            tlb_20_P1_MAT <= _GEN_2215;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_21_P0_PPN <= _GEN_966;
          end else begin
            tlb_21_P0_PPN <= _GEN_1992;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_21_P0_MAT <= _GEN_1030;
          end else begin
            tlb_21_P0_MAT <= _GEN_2056;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_21_P1_PPN <= _GEN_1126;
          end else begin
            tlb_21_P1_PPN <= _GEN_2152;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_21_P1_MAT <= _GEN_1190;
          end else begin
            tlb_21_P1_MAT <= _GEN_2216;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_22_P0_PPN <= _GEN_967;
          end else begin
            tlb_22_P0_PPN <= _GEN_1993;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_22_P0_MAT <= _GEN_1031;
          end else begin
            tlb_22_P0_MAT <= _GEN_2057;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_22_P1_PPN <= _GEN_1127;
          end else begin
            tlb_22_P1_PPN <= _GEN_2153;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_22_P1_MAT <= _GEN_1191;
          end else begin
            tlb_22_P1_MAT <= _GEN_2217;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_23_P0_PPN <= _GEN_968;
          end else begin
            tlb_23_P0_PPN <= _GEN_1994;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_23_P0_MAT <= _GEN_1032;
          end else begin
            tlb_23_P0_MAT <= _GEN_2058;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_23_P1_PPN <= _GEN_1128;
          end else begin
            tlb_23_P1_PPN <= _GEN_2154;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_23_P1_MAT <= _GEN_1192;
          end else begin
            tlb_23_P1_MAT <= _GEN_2218;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_24_P0_PPN <= _GEN_969;
          end else begin
            tlb_24_P0_PPN <= _GEN_1995;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_24_P0_MAT <= _GEN_1033;
          end else begin
            tlb_24_P0_MAT <= _GEN_2059;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_24_P1_PPN <= _GEN_1129;
          end else begin
            tlb_24_P1_PPN <= _GEN_2155;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_24_P1_MAT <= _GEN_1193;
          end else begin
            tlb_24_P1_MAT <= _GEN_2219;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_25_P0_PPN <= _GEN_970;
          end else begin
            tlb_25_P0_PPN <= _GEN_1996;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_25_P0_MAT <= _GEN_1034;
          end else begin
            tlb_25_P0_MAT <= _GEN_2060;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_25_P1_PPN <= _GEN_1130;
          end else begin
            tlb_25_P1_PPN <= _GEN_2156;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_25_P1_MAT <= _GEN_1194;
          end else begin
            tlb_25_P1_MAT <= _GEN_2220;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_26_P0_PPN <= _GEN_971;
          end else begin
            tlb_26_P0_PPN <= _GEN_1997;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_26_P0_MAT <= _GEN_1035;
          end else begin
            tlb_26_P0_MAT <= _GEN_2061;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_26_P1_PPN <= _GEN_1131;
          end else begin
            tlb_26_P1_PPN <= _GEN_2157;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_26_P1_MAT <= _GEN_1195;
          end else begin
            tlb_26_P1_MAT <= _GEN_2221;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_27_P0_PPN <= _GEN_972;
          end else begin
            tlb_27_P0_PPN <= _GEN_1998;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_27_P0_MAT <= _GEN_1036;
          end else begin
            tlb_27_P0_MAT <= _GEN_2062;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_27_P1_PPN <= _GEN_1132;
          end else begin
            tlb_27_P1_PPN <= _GEN_2158;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_27_P1_MAT <= _GEN_1196;
          end else begin
            tlb_27_P1_MAT <= _GEN_2222;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_28_P0_PPN <= _GEN_973;
          end else begin
            tlb_28_P0_PPN <= _GEN_1999;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_28_P0_MAT <= _GEN_1037;
          end else begin
            tlb_28_P0_MAT <= _GEN_2063;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_28_P1_PPN <= _GEN_1133;
          end else begin
            tlb_28_P1_PPN <= _GEN_2159;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_28_P1_MAT <= _GEN_1197;
          end else begin
            tlb_28_P1_MAT <= _GEN_2223;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_29_P0_PPN <= _GEN_974;
          end else begin
            tlb_29_P0_PPN <= _GEN_2000;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_29_P0_MAT <= _GEN_1038;
          end else begin
            tlb_29_P0_MAT <= _GEN_2064;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_29_P1_PPN <= _GEN_1134;
          end else begin
            tlb_29_P1_PPN <= _GEN_2160;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_29_P1_MAT <= _GEN_1198;
          end else begin
            tlb_29_P1_MAT <= _GEN_2224;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_30_P0_PPN <= _GEN_975;
          end else begin
            tlb_30_P0_PPN <= _GEN_2001;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_30_P0_MAT <= _GEN_1039;
          end else begin
            tlb_30_P0_MAT <= _GEN_2065;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_30_P1_PPN <= _GEN_1135;
          end else begin
            tlb_30_P1_PPN <= _GEN_2161;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_30_P1_MAT <= _GEN_1199;
          end else begin
            tlb_30_P1_MAT <= _GEN_2225;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_31_P0_PPN <= _GEN_976;
          end else begin
            tlb_31_P0_PPN <= _GEN_2002;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_31_P0_MAT <= _GEN_1040;
          end else begin
            tlb_31_P0_MAT <= _GEN_2066;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_31_P1_PPN <= _GEN_1136;
          end else begin
            tlb_31_P1_PPN <= _GEN_2162;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(_T_1443)) begin
        if (!(_T_1475)) begin
          if (_T_1476) begin
            tlb_31_P1_MAT <= _GEN_1200;
          end else begin
            tlb_31_P1_MAT <= _GEN_2226;
          end
        end
      end
    end
  end
endmodule
module SimpleLACoreWrapRAM(
  input         clock,
  input         reset,
  input         io_ipi,
  input  [7:0]  io_interrupt,
  output [31:0] io_debug_pc,
  output [3:0]  io_debug_wen,
  output [4:0]  io_debug_wnum,
  output [31:0] io_debug_wdata,
  output        io_inst_en,
  output [31:0] io_inst_addr,
  input  [31:0] io_inst_rdata,
  output        io_data_en,
  output [3:0]  io_data_wen,
  output [31:0] io_data_addr,
  output [31:0] io_data_wdata,
  input  [31:0] io_data_rdata
);
  wire  core_clock;
  wire  core_reset;
  wire  core_io_ipi;
  wire [7:0] core_io_interrupt;
  wire  core_io_inst_req_valid;
  wire [31:0] core_io_inst_req_bits_addr;
  wire  core_io_inst_resp_valid;
  wire [31:0] core_io_inst_resp_bits;
  wire  core_io_data_req_valid;
  wire [3:0] core_io_data_req_bits_wen;
  wire [31:0] core_io_data_req_bits_addr;
  wire [31:0] core_io_data_req_bits_wdata;
  wire  core_io_data_req_bits_cacop;
  wire  core_io_data_req_bits_preld;
  wire  core_io_data_resp_valid;
  wire [31:0] core_io_data_resp_bits;
  wire [31:0] core_io_debug_pc;
  wire [3:0] core_io_debug_wen;
  wire [4:0] core_io_debug_wnum;
  wire [31:0] core_io_debug_wdata;
  SimpleLACore core (
    .clock(core_clock),
    .reset(core_reset),
    .io_ipi(core_io_ipi),
    .io_interrupt(core_io_interrupt),
    .io_inst_req_valid(core_io_inst_req_valid),
    .io_inst_req_bits_addr(core_io_inst_req_bits_addr),
    .io_inst_resp_valid(core_io_inst_resp_valid),
    .io_inst_resp_bits(core_io_inst_resp_bits),
    .io_data_req_valid(core_io_data_req_valid),
    .io_data_req_bits_wen(core_io_data_req_bits_wen),
    .io_data_req_bits_addr(core_io_data_req_bits_addr),
    .io_data_req_bits_wdata(core_io_data_req_bits_wdata),
    .io_data_req_bits_cacop(core_io_data_req_bits_cacop),
    .io_data_req_bits_preld(core_io_data_req_bits_preld),
    .io_data_resp_valid(core_io_data_resp_valid),
    .io_data_resp_bits(core_io_data_resp_bits),
    .io_debug_pc(core_io_debug_pc),
    .io_debug_wen(core_io_debug_wen),
    .io_debug_wnum(core_io_debug_wnum),
    .io_debug_wdata(core_io_debug_wdata)
  );
  assign io_debug_pc = core_io_debug_pc;
  assign io_debug_wen = core_io_debug_wen;
  assign io_debug_wnum = core_io_debug_wnum;
  assign io_debug_wdata = core_io_debug_wdata;
  assign io_inst_en = core_io_inst_req_valid;
  assign io_inst_addr = core_io_inst_req_bits_addr;
  assign io_data_en = core_io_data_req_valid & ~core_io_data_req_bits_cacop & ~core_io_data_req_bits_preld;
  assign io_data_wen = core_io_data_req_bits_wen;
  assign io_data_addr = core_io_data_req_bits_addr;
  assign io_data_wdata = core_io_data_req_bits_wdata;
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_ipi = io_ipi;
  assign core_io_interrupt = io_interrupt;
  assign core_io_inst_resp_valid = core_io_inst_req_valid;
  assign core_io_inst_resp_bits = io_inst_rdata;
  assign core_io_data_resp_valid = core_io_data_req_valid;
  assign core_io_data_resp_bits = io_data_rdata;
endmodule
